pulp_write32(axi_m, 32'h44000000, 32'd0);
pulp_write32(axi_m, 32'h44000004, 32'd3);
pulp_write32(axi_m, 32'h44000008, 32'h80001928);
pulp_write32(axi_m, 32'h44001928, 32'h80000578);
pulp_write32(axi_m, 32'h4400192c, 32'h80000604);
pulp_write32(axi_m, 32'h44001930, 32'h80000690);
pulp_write32(axi_m, 32'h4400004c, 32'h00000000);
pulp_write32(axi_m, 32'h44000050, 32'h00000001);
pulp_write32(axi_m, 32'h44000054, 32'h00000002);
pulp_write32(axi_m, 32'h44000058, 32'h00000003);
pulp_write32(axi_m, 32'h4400005c, 32'h00000004);
pulp_write32(axi_m, 32'h44000060, 32'h00000005);
pulp_write32(axi_m, 32'h44000064, 32'h00000006);
pulp_write32(axi_m, 32'h44000068, 32'h00000007);
pulp_write32(axi_m, 32'h4400006c, 32'h00000008);
pulp_write32(axi_m, 32'h44000070, 32'h00000009);
pulp_write32(axi_m, 32'h44000074, 32'h0000000a);
pulp_write32(axi_m, 32'h44000078, 32'h0000000b);
pulp_write32(axi_m, 32'h4400007c, 32'h0000000c);
pulp_write32(axi_m, 32'h44000080, 32'h0000000d);
pulp_write32(axi_m, 32'h44000084, 32'h0000000e);
pulp_write32(axi_m, 32'h44000088, 32'h0000000f);

pulp_write32(axi_m, 32'h4400008c, 32'd1);
pulp_write32(axi_m, 32'h44000090, 32'd3);
pulp_write32(axi_m, 32'h44000094, 32'h80001938);
pulp_write32(axi_m, 32'h44001938, 32'h80000118);
pulp_write32(axi_m, 32'h4400193c, 32'h800003d4);
pulp_write32(axi_m, 32'h44001940, 32'h80000a64);
pulp_write32(axi_m, 32'h440000d8, 32'h00010000);
pulp_write32(axi_m, 32'h440000dc, 32'h00010001);
pulp_write32(axi_m, 32'h440000e0, 32'h00010002);
pulp_write32(axi_m, 32'h440000e4, 32'h00010003);
pulp_write32(axi_m, 32'h440000e8, 32'h00010004);
pulp_write32(axi_m, 32'h440000ec, 32'h00010005);
pulp_write32(axi_m, 32'h440000f0, 32'h00010006);
pulp_write32(axi_m, 32'h440000f4, 32'h00010007);
pulp_write32(axi_m, 32'h440000f8, 32'h00010008);
pulp_write32(axi_m, 32'h440000fc, 32'h00010009);
pulp_write32(axi_m, 32'h44000100, 32'h0001000a);
pulp_write32(axi_m, 32'h44000104, 32'h0001000b);
pulp_write32(axi_m, 32'h44000108, 32'h0001000c);
pulp_write32(axi_m, 32'h4400010c, 32'h0001000d);
pulp_write32(axi_m, 32'h44000110, 32'h0001000e);
pulp_write32(axi_m, 32'h44000114, 32'h0001000f);

pulp_write32(axi_m, 32'h44000118, 32'd2);
pulp_write32(axi_m, 32'h4400011c, 32'd2);
pulp_write32(axi_m, 32'h44000120, 32'h80001948);
pulp_write32(axi_m, 32'h44001948, 32'h800001a4);
pulp_write32(axi_m, 32'h4400194c, 32'h8000166c);
pulp_write32(axi_m, 32'h44000164, 32'h00020000);
pulp_write32(axi_m, 32'h44000168, 32'h00020001);
pulp_write32(axi_m, 32'h4400016c, 32'h00020002);
pulp_write32(axi_m, 32'h44000170, 32'h00020003);
pulp_write32(axi_m, 32'h44000174, 32'h00020004);
pulp_write32(axi_m, 32'h44000178, 32'h00020005);
pulp_write32(axi_m, 32'h4400017c, 32'h00020006);
pulp_write32(axi_m, 32'h44000180, 32'h00020007);
pulp_write32(axi_m, 32'h44000184, 32'h00020008);
pulp_write32(axi_m, 32'h44000188, 32'h00020009);
pulp_write32(axi_m, 32'h4400018c, 32'h0002000a);
pulp_write32(axi_m, 32'h44000190, 32'h0002000b);
pulp_write32(axi_m, 32'h44000194, 32'h0002000c);
pulp_write32(axi_m, 32'h44000198, 32'h0002000d);
pulp_write32(axi_m, 32'h4400019c, 32'h0002000e);
pulp_write32(axi_m, 32'h440001a0, 32'h0002000f);

pulp_write32(axi_m, 32'h440001a4, 32'd3);
pulp_write32(axi_m, 32'h440001a8, 32'd2);
pulp_write32(axi_m, 32'h440001ac, 32'h80001950);
pulp_write32(axi_m, 32'h44001950, 32'h80000230);
pulp_write32(axi_m, 32'h44001954, 32'h80000ec4);
pulp_write32(axi_m, 32'h440001f0, 32'h00030000);
pulp_write32(axi_m, 32'h440001f4, 32'h00030001);
pulp_write32(axi_m, 32'h440001f8, 32'h00030002);
pulp_write32(axi_m, 32'h440001fc, 32'h00030003);
pulp_write32(axi_m, 32'h44000200, 32'h00030004);
pulp_write32(axi_m, 32'h44000204, 32'h00030005);
pulp_write32(axi_m, 32'h44000208, 32'h00030006);
pulp_write32(axi_m, 32'h4400020c, 32'h00030007);
pulp_write32(axi_m, 32'h44000210, 32'h00030008);
pulp_write32(axi_m, 32'h44000214, 32'h00030009);
pulp_write32(axi_m, 32'h44000218, 32'h0003000a);
pulp_write32(axi_m, 32'h4400021c, 32'h0003000b);
pulp_write32(axi_m, 32'h44000220, 32'h0003000c);
pulp_write32(axi_m, 32'h44000224, 32'h0003000d);
pulp_write32(axi_m, 32'h44000228, 32'h0003000e);
pulp_write32(axi_m, 32'h4400022c, 32'h0003000f);

pulp_write32(axi_m, 32'h44000230, 32'd4);
pulp_write32(axi_m, 32'h44000234, 32'd2);
pulp_write32(axi_m, 32'h44000238, 32'h80001958);
pulp_write32(axi_m, 32'h44001958, 32'h800002bc);
pulp_write32(axi_m, 32'h4400195c, 32'h8000120c);
pulp_write32(axi_m, 32'h4400027c, 32'h00040000);
pulp_write32(axi_m, 32'h44000280, 32'h00040001);
pulp_write32(axi_m, 32'h44000284, 32'h00040002);
pulp_write32(axi_m, 32'h44000288, 32'h00040003);
pulp_write32(axi_m, 32'h4400028c, 32'h00040004);
pulp_write32(axi_m, 32'h44000290, 32'h00040005);
pulp_write32(axi_m, 32'h44000294, 32'h00040006);
pulp_write32(axi_m, 32'h44000298, 32'h00040007);
pulp_write32(axi_m, 32'h4400029c, 32'h00040008);
pulp_write32(axi_m, 32'h440002a0, 32'h00040009);
pulp_write32(axi_m, 32'h440002a4, 32'h0004000a);
pulp_write32(axi_m, 32'h440002a8, 32'h0004000b);
pulp_write32(axi_m, 32'h440002ac, 32'h0004000c);
pulp_write32(axi_m, 32'h440002b0, 32'h0004000d);
pulp_write32(axi_m, 32'h440002b4, 32'h0004000e);
pulp_write32(axi_m, 32'h440002b8, 32'h0004000f);

pulp_write32(axi_m, 32'h440002bc, 32'd5);
pulp_write32(axi_m, 32'h440002c0, 32'd2);
pulp_write32(axi_m, 32'h440002c4, 32'h80001960);
pulp_write32(axi_m, 32'h44001960, 32'h80000348);
pulp_write32(axi_m, 32'h44001964, 32'h8000189c);
pulp_write32(axi_m, 32'h44000308, 32'h00050000);
pulp_write32(axi_m, 32'h4400030c, 32'h00050001);
pulp_write32(axi_m, 32'h44000310, 32'h00050002);
pulp_write32(axi_m, 32'h44000314, 32'h00050003);
pulp_write32(axi_m, 32'h44000318, 32'h00050004);
pulp_write32(axi_m, 32'h4400031c, 32'h00050005);
pulp_write32(axi_m, 32'h44000320, 32'h00050006);
pulp_write32(axi_m, 32'h44000324, 32'h00050007);
pulp_write32(axi_m, 32'h44000328, 32'h00050008);
pulp_write32(axi_m, 32'h4400032c, 32'h00050009);
pulp_write32(axi_m, 32'h44000330, 32'h0005000a);
pulp_write32(axi_m, 32'h44000334, 32'h0005000b);
pulp_write32(axi_m, 32'h44000338, 32'h0005000c);
pulp_write32(axi_m, 32'h4400033c, 32'h0005000d);
pulp_write32(axi_m, 32'h44000340, 32'h0005000e);
pulp_write32(axi_m, 32'h44000344, 32'h0005000f);

pulp_write32(axi_m, 32'h44000348, 32'd6);
pulp_write32(axi_m, 32'h4400034c, 32'd2);
pulp_write32(axi_m, 32'h44000350, 32'h80001968);
pulp_write32(axi_m, 32'h44001968, 32'h800004ec);
pulp_write32(axi_m, 32'h4400196c, 32'h80000fdc);
pulp_write32(axi_m, 32'h44000394, 32'h00060000);
pulp_write32(axi_m, 32'h44000398, 32'h00060001);
pulp_write32(axi_m, 32'h4400039c, 32'h00060002);
pulp_write32(axi_m, 32'h440003a0, 32'h00060003);
pulp_write32(axi_m, 32'h440003a4, 32'h00060004);
pulp_write32(axi_m, 32'h440003a8, 32'h00060005);
pulp_write32(axi_m, 32'h440003ac, 32'h00060006);
pulp_write32(axi_m, 32'h440003b0, 32'h00060007);
pulp_write32(axi_m, 32'h440003b4, 32'h00060008);
pulp_write32(axi_m, 32'h440003b8, 32'h00060009);
pulp_write32(axi_m, 32'h440003bc, 32'h0006000a);
pulp_write32(axi_m, 32'h440003c0, 32'h0006000b);
pulp_write32(axi_m, 32'h440003c4, 32'h0006000c);
pulp_write32(axi_m, 32'h440003c8, 32'h0006000d);
pulp_write32(axi_m, 32'h440003cc, 32'h0006000e);
pulp_write32(axi_m, 32'h440003d0, 32'h0006000f);

pulp_write32(axi_m, 32'h440003d4, 32'd7);
pulp_write32(axi_m, 32'h440003d8, 32'd2);
pulp_write32(axi_m, 32'h440003dc, 32'h80001970);
pulp_write32(axi_m, 32'h44001970, 32'h80000460);
pulp_write32(axi_m, 32'h44001974, 32'h80000b7c);
pulp_write32(axi_m, 32'h44000420, 32'h00070000);
pulp_write32(axi_m, 32'h44000424, 32'h00070001);
pulp_write32(axi_m, 32'h44000428, 32'h00070002);
pulp_write32(axi_m, 32'h4400042c, 32'h00070003);
pulp_write32(axi_m, 32'h44000430, 32'h00070004);
pulp_write32(axi_m, 32'h44000434, 32'h00070005);
pulp_write32(axi_m, 32'h44000438, 32'h00070006);
pulp_write32(axi_m, 32'h4400043c, 32'h00070007);
pulp_write32(axi_m, 32'h44000440, 32'h00070008);
pulp_write32(axi_m, 32'h44000444, 32'h00070009);
pulp_write32(axi_m, 32'h44000448, 32'h0007000a);
pulp_write32(axi_m, 32'h4400044c, 32'h0007000b);
pulp_write32(axi_m, 32'h44000450, 32'h0007000c);
pulp_write32(axi_m, 32'h44000454, 32'h0007000d);
pulp_write32(axi_m, 32'h44000458, 32'h0007000e);
pulp_write32(axi_m, 32'h4400045c, 32'h0007000f);

pulp_write32(axi_m, 32'h44000460, 32'd8);
pulp_write32(axi_m, 32'h44000464, 32'd2);
pulp_write32(axi_m, 32'h44000468, 32'h80001978);
pulp_write32(axi_m, 32'h44001978, 32'h800004ec);
pulp_write32(axi_m, 32'h4400197c, 32'h80000c08);
pulp_write32(axi_m, 32'h440004ac, 32'h00080000);
pulp_write32(axi_m, 32'h440004b0, 32'h00080001);
pulp_write32(axi_m, 32'h440004b4, 32'h00080002);
pulp_write32(axi_m, 32'h440004b8, 32'h00080003);
pulp_write32(axi_m, 32'h440004bc, 32'h00080004);
pulp_write32(axi_m, 32'h440004c0, 32'h00080005);
pulp_write32(axi_m, 32'h440004c4, 32'h00080006);
pulp_write32(axi_m, 32'h440004c8, 32'h00080007);
pulp_write32(axi_m, 32'h440004cc, 32'h00080008);
pulp_write32(axi_m, 32'h440004d0, 32'h00080009);
pulp_write32(axi_m, 32'h440004d4, 32'h0008000a);
pulp_write32(axi_m, 32'h440004d8, 32'h0008000b);
pulp_write32(axi_m, 32'h440004dc, 32'h0008000c);
pulp_write32(axi_m, 32'h440004e0, 32'h0008000d);
pulp_write32(axi_m, 32'h440004e4, 32'h0008000e);
pulp_write32(axi_m, 32'h440004e8, 32'h0008000f);

pulp_write32(axi_m, 32'h440004ec, 32'd9);
pulp_write32(axi_m, 32'h440004f0, 32'd1);
pulp_write32(axi_m, 32'h440004f4, 32'h80001980);
pulp_write32(axi_m, 32'h44001980, 32'h80000d20);
pulp_write32(axi_m, 32'h44000538, 32'h00090000);
pulp_write32(axi_m, 32'h4400053c, 32'h00090001);
pulp_write32(axi_m, 32'h44000540, 32'h00090002);
pulp_write32(axi_m, 32'h44000544, 32'h00090003);
pulp_write32(axi_m, 32'h44000548, 32'h00090004);
pulp_write32(axi_m, 32'h4400054c, 32'h00090005);
pulp_write32(axi_m, 32'h44000550, 32'h00090006);
pulp_write32(axi_m, 32'h44000554, 32'h00090007);
pulp_write32(axi_m, 32'h44000558, 32'h00090008);
pulp_write32(axi_m, 32'h4400055c, 32'h00090009);
pulp_write32(axi_m, 32'h44000560, 32'h0009000a);
pulp_write32(axi_m, 32'h44000564, 32'h0009000b);
pulp_write32(axi_m, 32'h44000568, 32'h0009000c);
pulp_write32(axi_m, 32'h4400056c, 32'h0009000d);
pulp_write32(axi_m, 32'h44000570, 32'h0009000e);
pulp_write32(axi_m, 32'h44000574, 32'h0009000f);

pulp_write32(axi_m, 32'h44000578, 32'd10);
pulp_write32(axi_m, 32'h4400057c, 32'd2);
pulp_write32(axi_m, 32'h44000580, 32'h80001988);
pulp_write32(axi_m, 32'h44001988, 32'h8000071c);
pulp_write32(axi_m, 32'h4400198c, 32'h800007a8);
pulp_write32(axi_m, 32'h440005c4, 32'h000a0000);
pulp_write32(axi_m, 32'h440005c8, 32'h000a0001);
pulp_write32(axi_m, 32'h440005cc, 32'h000a0002);
pulp_write32(axi_m, 32'h440005d0, 32'h000a0003);
pulp_write32(axi_m, 32'h440005d4, 32'h000a0004);
pulp_write32(axi_m, 32'h440005d8, 32'h000a0005);
pulp_write32(axi_m, 32'h440005dc, 32'h000a0006);
pulp_write32(axi_m, 32'h440005e0, 32'h000a0007);
pulp_write32(axi_m, 32'h440005e4, 32'h000a0008);
pulp_write32(axi_m, 32'h440005e8, 32'h000a0009);
pulp_write32(axi_m, 32'h440005ec, 32'h000a000a);
pulp_write32(axi_m, 32'h440005f0, 32'h000a000b);
pulp_write32(axi_m, 32'h440005f4, 32'h000a000c);
pulp_write32(axi_m, 32'h440005f8, 32'h000a000d);
pulp_write32(axi_m, 32'h440005fc, 32'h000a000e);
pulp_write32(axi_m, 32'h44000600, 32'h000a000f);

pulp_write32(axi_m, 32'h44000604, 32'd11);
pulp_write32(axi_m, 32'h44000608, 32'd2);
pulp_write32(axi_m, 32'h4400060c, 32'h80001990);
pulp_write32(axi_m, 32'h44001990, 32'h80000e38);
pulp_write32(axi_m, 32'h44001994, 32'h80000f50);
pulp_write32(axi_m, 32'h44000650, 32'h000b0000);
pulp_write32(axi_m, 32'h44000654, 32'h000b0001);
pulp_write32(axi_m, 32'h44000658, 32'h000b0002);
pulp_write32(axi_m, 32'h4400065c, 32'h000b0003);
pulp_write32(axi_m, 32'h44000660, 32'h000b0004);
pulp_write32(axi_m, 32'h44000664, 32'h000b0005);
pulp_write32(axi_m, 32'h44000668, 32'h000b0006);
pulp_write32(axi_m, 32'h4400066c, 32'h000b0007);
pulp_write32(axi_m, 32'h44000670, 32'h000b0008);
pulp_write32(axi_m, 32'h44000674, 32'h000b0009);
pulp_write32(axi_m, 32'h44000678, 32'h000b000a);
pulp_write32(axi_m, 32'h4400067c, 32'h000b000b);
pulp_write32(axi_m, 32'h44000680, 32'h000b000c);
pulp_write32(axi_m, 32'h44000684, 32'h000b000d);
pulp_write32(axi_m, 32'h44000688, 32'h000b000e);
pulp_write32(axi_m, 32'h4400068c, 32'h000b000f);

pulp_write32(axi_m, 32'h44000690, 32'd12);
pulp_write32(axi_m, 32'h44000694, 32'd2);
pulp_write32(axi_m, 32'h44000698, 32'h80001998);
pulp_write32(axi_m, 32'h44001998, 32'h80001068);
pulp_write32(axi_m, 32'h4400199c, 32'h800010f4);
pulp_write32(axi_m, 32'h440006dc, 32'h000c0000);
pulp_write32(axi_m, 32'h440006e0, 32'h000c0001);
pulp_write32(axi_m, 32'h440006e4, 32'h000c0002);
pulp_write32(axi_m, 32'h440006e8, 32'h000c0003);
pulp_write32(axi_m, 32'h440006ec, 32'h000c0004);
pulp_write32(axi_m, 32'h440006f0, 32'h000c0005);
pulp_write32(axi_m, 32'h440006f4, 32'h000c0006);
pulp_write32(axi_m, 32'h440006f8, 32'h000c0007);
pulp_write32(axi_m, 32'h440006fc, 32'h000c0008);
pulp_write32(axi_m, 32'h44000700, 32'h000c0009);
pulp_write32(axi_m, 32'h44000704, 32'h000c000a);
pulp_write32(axi_m, 32'h44000708, 32'h000c000b);
pulp_write32(axi_m, 32'h4400070c, 32'h000c000c);
pulp_write32(axi_m, 32'h44000710, 32'h000c000d);
pulp_write32(axi_m, 32'h44000714, 32'h000c000e);
pulp_write32(axi_m, 32'h44000718, 32'h000c000f);

pulp_write32(axi_m, 32'h4400071c, 32'd13);
pulp_write32(axi_m, 32'h44000720, 32'd2);
pulp_write32(axi_m, 32'h44000724, 32'h800019a0);
pulp_write32(axi_m, 32'h440019a0, 32'h80000834);
pulp_write32(axi_m, 32'h440019a4, 32'h80000b7c);
pulp_write32(axi_m, 32'h44000768, 32'h000d0000);
pulp_write32(axi_m, 32'h4400076c, 32'h000d0001);
pulp_write32(axi_m, 32'h44000770, 32'h000d0002);
pulp_write32(axi_m, 32'h44000774, 32'h000d0003);
pulp_write32(axi_m, 32'h44000778, 32'h000d0004);
pulp_write32(axi_m, 32'h4400077c, 32'h000d0005);
pulp_write32(axi_m, 32'h44000780, 32'h000d0006);
pulp_write32(axi_m, 32'h44000784, 32'h000d0007);
pulp_write32(axi_m, 32'h44000788, 32'h000d0008);
pulp_write32(axi_m, 32'h4400078c, 32'h000d0009);
pulp_write32(axi_m, 32'h44000790, 32'h000d000a);
pulp_write32(axi_m, 32'h44000794, 32'h000d000b);
pulp_write32(axi_m, 32'h44000798, 32'h000d000c);
pulp_write32(axi_m, 32'h4400079c, 32'h000d000d);
pulp_write32(axi_m, 32'h440007a0, 32'h000d000e);
pulp_write32(axi_m, 32'h440007a4, 32'h000d000f);

pulp_write32(axi_m, 32'h440007a8, 32'd14);
pulp_write32(axi_m, 32'h440007ac, 32'd2);
pulp_write32(axi_m, 32'h440007b0, 32'h800019a8);
pulp_write32(axi_m, 32'h440019a8, 32'h80000834);
pulp_write32(axi_m, 32'h440019ac, 32'h800009d8);
pulp_write32(axi_m, 32'h440007f4, 32'h000e0000);
pulp_write32(axi_m, 32'h440007f8, 32'h000e0001);
pulp_write32(axi_m, 32'h440007fc, 32'h000e0002);
pulp_write32(axi_m, 32'h44000800, 32'h000e0003);
pulp_write32(axi_m, 32'h44000804, 32'h000e0004);
pulp_write32(axi_m, 32'h44000808, 32'h000e0005);
pulp_write32(axi_m, 32'h4400080c, 32'h000e0006);
pulp_write32(axi_m, 32'h44000810, 32'h000e0007);
pulp_write32(axi_m, 32'h44000814, 32'h000e0008);
pulp_write32(axi_m, 32'h44000818, 32'h000e0009);
pulp_write32(axi_m, 32'h4400081c, 32'h000e000a);
pulp_write32(axi_m, 32'h44000820, 32'h000e000b);
pulp_write32(axi_m, 32'h44000824, 32'h000e000c);
pulp_write32(axi_m, 32'h44000828, 32'h000e000d);
pulp_write32(axi_m, 32'h4400082c, 32'h000e000e);
pulp_write32(axi_m, 32'h44000830, 32'h000e000f);

pulp_write32(axi_m, 32'h44000834, 32'd15);
pulp_write32(axi_m, 32'h44000838, 32'd1);
pulp_write32(axi_m, 32'h4400083c, 32'h800019b0);
pulp_write32(axi_m, 32'h440019b0, 32'h800008c0);
pulp_write32(axi_m, 32'h44000880, 32'h000f0000);
pulp_write32(axi_m, 32'h44000884, 32'h000f0001);
pulp_write32(axi_m, 32'h44000888, 32'h000f0002);
pulp_write32(axi_m, 32'h4400088c, 32'h000f0003);
pulp_write32(axi_m, 32'h44000890, 32'h000f0004);
pulp_write32(axi_m, 32'h44000894, 32'h000f0005);
pulp_write32(axi_m, 32'h44000898, 32'h000f0006);
pulp_write32(axi_m, 32'h4400089c, 32'h000f0007);
pulp_write32(axi_m, 32'h440008a0, 32'h000f0008);
pulp_write32(axi_m, 32'h440008a4, 32'h000f0009);
pulp_write32(axi_m, 32'h440008a8, 32'h000f000a);
pulp_write32(axi_m, 32'h440008ac, 32'h000f000b);
pulp_write32(axi_m, 32'h440008b0, 32'h000f000c);
pulp_write32(axi_m, 32'h440008b4, 32'h000f000d);
pulp_write32(axi_m, 32'h440008b8, 32'h000f000e);
pulp_write32(axi_m, 32'h440008bc, 32'h000f000f);

pulp_write32(axi_m, 32'h440008c0, 32'd16);
pulp_write32(axi_m, 32'h440008c4, 32'd2);
pulp_write32(axi_m, 32'h440008c8, 32'h800019b8);
pulp_write32(axi_m, 32'h440019b8, 32'h8000094c);
pulp_write32(axi_m, 32'h440019bc, 32'h80000af0);
pulp_write32(axi_m, 32'h4400090c, 32'h00100000);
pulp_write32(axi_m, 32'h44000910, 32'h00100001);
pulp_write32(axi_m, 32'h44000914, 32'h00100002);
pulp_write32(axi_m, 32'h44000918, 32'h00100003);
pulp_write32(axi_m, 32'h4400091c, 32'h00100004);
pulp_write32(axi_m, 32'h44000920, 32'h00100005);
pulp_write32(axi_m, 32'h44000924, 32'h00100006);
pulp_write32(axi_m, 32'h44000928, 32'h00100007);
pulp_write32(axi_m, 32'h4400092c, 32'h00100008);
pulp_write32(axi_m, 32'h44000930, 32'h00100009);
pulp_write32(axi_m, 32'h44000934, 32'h0010000a);
pulp_write32(axi_m, 32'h44000938, 32'h0010000b);
pulp_write32(axi_m, 32'h4400093c, 32'h0010000c);
pulp_write32(axi_m, 32'h44000940, 32'h0010000d);
pulp_write32(axi_m, 32'h44000944, 32'h0010000e);
pulp_write32(axi_m, 32'h44000948, 32'h0010000f);

pulp_write32(axi_m, 32'h4400094c, 32'd17);
pulp_write32(axi_m, 32'h44000950, 32'd2);
pulp_write32(axi_m, 32'h44000954, 32'h800019c0);
pulp_write32(axi_m, 32'h440019c0, 32'h800009d8);
pulp_write32(axi_m, 32'h440019c4, 32'h80000c94);
pulp_write32(axi_m, 32'h44000998, 32'h00110000);
pulp_write32(axi_m, 32'h4400099c, 32'h00110001);
pulp_write32(axi_m, 32'h440009a0, 32'h00110002);
pulp_write32(axi_m, 32'h440009a4, 32'h00110003);
pulp_write32(axi_m, 32'h440009a8, 32'h00110004);
pulp_write32(axi_m, 32'h440009ac, 32'h00110005);
pulp_write32(axi_m, 32'h440009b0, 32'h00110006);
pulp_write32(axi_m, 32'h440009b4, 32'h00110007);
pulp_write32(axi_m, 32'h440009b8, 32'h00110008);
pulp_write32(axi_m, 32'h440009bc, 32'h00110009);
pulp_write32(axi_m, 32'h440009c0, 32'h0011000a);
pulp_write32(axi_m, 32'h440009c4, 32'h0011000b);
pulp_write32(axi_m, 32'h440009c8, 32'h0011000c);
pulp_write32(axi_m, 32'h440009cc, 32'h0011000d);
pulp_write32(axi_m, 32'h440009d0, 32'h0011000e);
pulp_write32(axi_m, 32'h440009d4, 32'h0011000f);

pulp_write32(axi_m, 32'h440009d8, 32'd18);
pulp_write32(axi_m, 32'h440009dc, 32'd1);
pulp_write32(axi_m, 32'h440009e0, 32'h800019c8);
pulp_write32(axi_m, 32'h440019c8, 32'h80000d20);
pulp_write32(axi_m, 32'h44000a24, 32'h00120000);
pulp_write32(axi_m, 32'h44000a28, 32'h00120001);
pulp_write32(axi_m, 32'h44000a2c, 32'h00120002);
pulp_write32(axi_m, 32'h44000a30, 32'h00120003);
pulp_write32(axi_m, 32'h44000a34, 32'h00120004);
pulp_write32(axi_m, 32'h44000a38, 32'h00120005);
pulp_write32(axi_m, 32'h44000a3c, 32'h00120006);
pulp_write32(axi_m, 32'h44000a40, 32'h00120007);
pulp_write32(axi_m, 32'h44000a44, 32'h00120008);
pulp_write32(axi_m, 32'h44000a48, 32'h00120009);
pulp_write32(axi_m, 32'h44000a4c, 32'h0012000a);
pulp_write32(axi_m, 32'h44000a50, 32'h0012000b);
pulp_write32(axi_m, 32'h44000a54, 32'h0012000c);
pulp_write32(axi_m, 32'h44000a58, 32'h0012000d);
pulp_write32(axi_m, 32'h44000a5c, 32'h0012000e);
pulp_write32(axi_m, 32'h44000a60, 32'h0012000f);

pulp_write32(axi_m, 32'h44000a64, 32'd19);
pulp_write32(axi_m, 32'h44000a68, 32'd2);
pulp_write32(axi_m, 32'h44000a6c, 32'h800019d0);
pulp_write32(axi_m, 32'h440019d0, 32'h80000dac);
pulp_write32(axi_m, 32'h440019d4, 32'h800015e0);
pulp_write32(axi_m, 32'h44000ab0, 32'h00130000);
pulp_write32(axi_m, 32'h44000ab4, 32'h00130001);
pulp_write32(axi_m, 32'h44000ab8, 32'h00130002);
pulp_write32(axi_m, 32'h44000abc, 32'h00130003);
pulp_write32(axi_m, 32'h44000ac0, 32'h00130004);
pulp_write32(axi_m, 32'h44000ac4, 32'h00130005);
pulp_write32(axi_m, 32'h44000ac8, 32'h00130006);
pulp_write32(axi_m, 32'h44000acc, 32'h00130007);
pulp_write32(axi_m, 32'h44000ad0, 32'h00130008);
pulp_write32(axi_m, 32'h44000ad4, 32'h00130009);
pulp_write32(axi_m, 32'h44000ad8, 32'h0013000a);
pulp_write32(axi_m, 32'h44000adc, 32'h0013000b);
pulp_write32(axi_m, 32'h44000ae0, 32'h0013000c);
pulp_write32(axi_m, 32'h44000ae4, 32'h0013000d);
pulp_write32(axi_m, 32'h44000ae8, 32'h0013000e);
pulp_write32(axi_m, 32'h44000aec, 32'h0013000f);

pulp_write32(axi_m, 32'h44000af0, 32'd20);
pulp_write32(axi_m, 32'h44000af4, 32'd2);
pulp_write32(axi_m, 32'h44000af8, 32'h800019d8);
pulp_write32(axi_m, 32'h440019d8, 32'h80000b7c);
pulp_write32(axi_m, 32'h440019dc, 32'h80000c08);
pulp_write32(axi_m, 32'h44000b3c, 32'h00140000);
pulp_write32(axi_m, 32'h44000b40, 32'h00140001);
pulp_write32(axi_m, 32'h44000b44, 32'h00140002);
pulp_write32(axi_m, 32'h44000b48, 32'h00140003);
pulp_write32(axi_m, 32'h44000b4c, 32'h00140004);
pulp_write32(axi_m, 32'h44000b50, 32'h00140005);
pulp_write32(axi_m, 32'h44000b54, 32'h00140006);
pulp_write32(axi_m, 32'h44000b58, 32'h00140007);
pulp_write32(axi_m, 32'h44000b5c, 32'h00140008);
pulp_write32(axi_m, 32'h44000b60, 32'h00140009);
pulp_write32(axi_m, 32'h44000b64, 32'h0014000a);
pulp_write32(axi_m, 32'h44000b68, 32'h0014000b);
pulp_write32(axi_m, 32'h44000b6c, 32'h0014000c);
pulp_write32(axi_m, 32'h44000b70, 32'h0014000d);
pulp_write32(axi_m, 32'h44000b74, 32'h0014000e);
pulp_write32(axi_m, 32'h44000b78, 32'h0014000f);

pulp_write32(axi_m, 32'h44000b7c, 32'd21);
pulp_write32(axi_m, 32'h44000b80, 32'd0);
pulp_write32(axi_m, 32'h44000bc8, 32'h00150000);
pulp_write32(axi_m, 32'h44000bcc, 32'h00150001);
pulp_write32(axi_m, 32'h44000bd0, 32'h00150002);
pulp_write32(axi_m, 32'h44000bd4, 32'h00150003);
pulp_write32(axi_m, 32'h44000bd8, 32'h00150004);
pulp_write32(axi_m, 32'h44000bdc, 32'h00150005);
pulp_write32(axi_m, 32'h44000be0, 32'h00150006);
pulp_write32(axi_m, 32'h44000be4, 32'h00150007);
pulp_write32(axi_m, 32'h44000be8, 32'h00150008);
pulp_write32(axi_m, 32'h44000bec, 32'h00150009);
pulp_write32(axi_m, 32'h44000bf0, 32'h0015000a);
pulp_write32(axi_m, 32'h44000bf4, 32'h0015000b);
pulp_write32(axi_m, 32'h44000bf8, 32'h0015000c);
pulp_write32(axi_m, 32'h44000bfc, 32'h0015000d);
pulp_write32(axi_m, 32'h44000c00, 32'h0015000e);
pulp_write32(axi_m, 32'h44000c04, 32'h0015000f);

pulp_write32(axi_m, 32'h44000c08, 32'd22);
pulp_write32(axi_m, 32'h44000c0c, 32'd1);
pulp_write32(axi_m, 32'h44000c10, 32'h800019e0);
pulp_write32(axi_m, 32'h440019e0, 32'h80000c94);
pulp_write32(axi_m, 32'h44000c54, 32'h00160000);
pulp_write32(axi_m, 32'h44000c58, 32'h00160001);
pulp_write32(axi_m, 32'h44000c5c, 32'h00160002);
pulp_write32(axi_m, 32'h44000c60, 32'h00160003);
pulp_write32(axi_m, 32'h44000c64, 32'h00160004);
pulp_write32(axi_m, 32'h44000c68, 32'h00160005);
pulp_write32(axi_m, 32'h44000c6c, 32'h00160006);
pulp_write32(axi_m, 32'h44000c70, 32'h00160007);
pulp_write32(axi_m, 32'h44000c74, 32'h00160008);
pulp_write32(axi_m, 32'h44000c78, 32'h00160009);
pulp_write32(axi_m, 32'h44000c7c, 32'h0016000a);
pulp_write32(axi_m, 32'h44000c80, 32'h0016000b);
pulp_write32(axi_m, 32'h44000c84, 32'h0016000c);
pulp_write32(axi_m, 32'h44000c88, 32'h0016000d);
pulp_write32(axi_m, 32'h44000c8c, 32'h0016000e);
pulp_write32(axi_m, 32'h44000c90, 32'h0016000f);

pulp_write32(axi_m, 32'h44000c94, 32'd23);
pulp_write32(axi_m, 32'h44000c98, 32'd1);
pulp_write32(axi_m, 32'h44000c9c, 32'h800019e8);
pulp_write32(axi_m, 32'h440019e8, 32'h80000d20);
pulp_write32(axi_m, 32'h44000ce0, 32'h00170000);
pulp_write32(axi_m, 32'h44000ce4, 32'h00170001);
pulp_write32(axi_m, 32'h44000ce8, 32'h00170002);
pulp_write32(axi_m, 32'h44000cec, 32'h00170003);
pulp_write32(axi_m, 32'h44000cf0, 32'h00170004);
pulp_write32(axi_m, 32'h44000cf4, 32'h00170005);
pulp_write32(axi_m, 32'h44000cf8, 32'h00170006);
pulp_write32(axi_m, 32'h44000cfc, 32'h00170007);
pulp_write32(axi_m, 32'h44000d00, 32'h00170008);
pulp_write32(axi_m, 32'h44000d04, 32'h00170009);
pulp_write32(axi_m, 32'h44000d08, 32'h0017000a);
pulp_write32(axi_m, 32'h44000d0c, 32'h0017000b);
pulp_write32(axi_m, 32'h44000d10, 32'h0017000c);
pulp_write32(axi_m, 32'h44000d14, 32'h0017000d);
pulp_write32(axi_m, 32'h44000d18, 32'h0017000e);
pulp_write32(axi_m, 32'h44000d1c, 32'h0017000f);

pulp_write32(axi_m, 32'h44000d20, 32'd24);
pulp_write32(axi_m, 32'h44000d24, 32'd0);
pulp_write32(axi_m, 32'h44000d6c, 32'h00180000);
pulp_write32(axi_m, 32'h44000d70, 32'h00180001);
pulp_write32(axi_m, 32'h44000d74, 32'h00180002);
pulp_write32(axi_m, 32'h44000d78, 32'h00180003);
pulp_write32(axi_m, 32'h44000d7c, 32'h00180004);
pulp_write32(axi_m, 32'h44000d80, 32'h00180005);
pulp_write32(axi_m, 32'h44000d84, 32'h00180006);
pulp_write32(axi_m, 32'h44000d88, 32'h00180007);
pulp_write32(axi_m, 32'h44000d8c, 32'h00180008);
pulp_write32(axi_m, 32'h44000d90, 32'h00180009);
pulp_write32(axi_m, 32'h44000d94, 32'h0018000a);
pulp_write32(axi_m, 32'h44000d98, 32'h0018000b);
pulp_write32(axi_m, 32'h44000d9c, 32'h0018000c);
pulp_write32(axi_m, 32'h44000da0, 32'h0018000d);
pulp_write32(axi_m, 32'h44000da4, 32'h0018000e);
pulp_write32(axi_m, 32'h44000da8, 32'h0018000f);

pulp_write32(axi_m, 32'h44000dac, 32'd25);
pulp_write32(axi_m, 32'h44000db0, 32'd2);
pulp_write32(axi_m, 32'h44000db4, 32'h800019f0);
pulp_write32(axi_m, 32'h440019f0, 32'h80000e38);
pulp_write32(axi_m, 32'h440019f4, 32'h800014c8);
pulp_write32(axi_m, 32'h44000df8, 32'h00190000);
pulp_write32(axi_m, 32'h44000dfc, 32'h00190001);
pulp_write32(axi_m, 32'h44000e00, 32'h00190002);
pulp_write32(axi_m, 32'h44000e04, 32'h00190003);
pulp_write32(axi_m, 32'h44000e08, 32'h00190004);
pulp_write32(axi_m, 32'h44000e0c, 32'h00190005);
pulp_write32(axi_m, 32'h44000e10, 32'h00190006);
pulp_write32(axi_m, 32'h44000e14, 32'h00190007);
pulp_write32(axi_m, 32'h44000e18, 32'h00190008);
pulp_write32(axi_m, 32'h44000e1c, 32'h00190009);
pulp_write32(axi_m, 32'h44000e20, 32'h0019000a);
pulp_write32(axi_m, 32'h44000e24, 32'h0019000b);
pulp_write32(axi_m, 32'h44000e28, 32'h0019000c);
pulp_write32(axi_m, 32'h44000e2c, 32'h0019000d);
pulp_write32(axi_m, 32'h44000e30, 32'h0019000e);
pulp_write32(axi_m, 32'h44000e34, 32'h0019000f);

pulp_write32(axi_m, 32'h44000e38, 32'd26);
pulp_write32(axi_m, 32'h44000e3c, 32'd1);
pulp_write32(axi_m, 32'h44000e40, 32'h800019f8);
pulp_write32(axi_m, 32'h440019f8, 32'h80001298);
pulp_write32(axi_m, 32'h44000e84, 32'h001a0000);
pulp_write32(axi_m, 32'h44000e88, 32'h001a0001);
pulp_write32(axi_m, 32'h44000e8c, 32'h001a0002);
pulp_write32(axi_m, 32'h44000e90, 32'h001a0003);
pulp_write32(axi_m, 32'h44000e94, 32'h001a0004);
pulp_write32(axi_m, 32'h44000e98, 32'h001a0005);
pulp_write32(axi_m, 32'h44000e9c, 32'h001a0006);
pulp_write32(axi_m, 32'h44000ea0, 32'h001a0007);
pulp_write32(axi_m, 32'h44000ea4, 32'h001a0008);
pulp_write32(axi_m, 32'h44000ea8, 32'h001a0009);
pulp_write32(axi_m, 32'h44000eac, 32'h001a000a);
pulp_write32(axi_m, 32'h44000eb0, 32'h001a000b);
pulp_write32(axi_m, 32'h44000eb4, 32'h001a000c);
pulp_write32(axi_m, 32'h44000eb8, 32'h001a000d);
pulp_write32(axi_m, 32'h44000ebc, 32'h001a000e);
pulp_write32(axi_m, 32'h44000ec0, 32'h001a000f);

pulp_write32(axi_m, 32'h44000ec4, 32'd27);
pulp_write32(axi_m, 32'h44000ec8, 32'd2);
pulp_write32(axi_m, 32'h44000ecc, 32'h80001a00);
pulp_write32(axi_m, 32'h44001a00, 32'h80000f50);
pulp_write32(axi_m, 32'h44001a04, 32'h80001554);
pulp_write32(axi_m, 32'h44000f10, 32'h001b0000);
pulp_write32(axi_m, 32'h44000f14, 32'h001b0001);
pulp_write32(axi_m, 32'h44000f18, 32'h001b0002);
pulp_write32(axi_m, 32'h44000f1c, 32'h001b0003);
pulp_write32(axi_m, 32'h44000f20, 32'h001b0004);
pulp_write32(axi_m, 32'h44000f24, 32'h001b0005);
pulp_write32(axi_m, 32'h44000f28, 32'h001b0006);
pulp_write32(axi_m, 32'h44000f2c, 32'h001b0007);
pulp_write32(axi_m, 32'h44000f30, 32'h001b0008);
pulp_write32(axi_m, 32'h44000f34, 32'h001b0009);
pulp_write32(axi_m, 32'h44000f38, 32'h001b000a);
pulp_write32(axi_m, 32'h44000f3c, 32'h001b000b);
pulp_write32(axi_m, 32'h44000f40, 32'h001b000c);
pulp_write32(axi_m, 32'h44000f44, 32'h001b000d);
pulp_write32(axi_m, 32'h44000f48, 32'h001b000e);
pulp_write32(axi_m, 32'h44000f4c, 32'h001b000f);

pulp_write32(axi_m, 32'h44000f50, 32'd28);
pulp_write32(axi_m, 32'h44000f54, 32'd1);
pulp_write32(axi_m, 32'h44000f58, 32'h80001a08);
pulp_write32(axi_m, 32'h44001a08, 32'h80001298);
pulp_write32(axi_m, 32'h44000f9c, 32'h001c0000);
pulp_write32(axi_m, 32'h44000fa0, 32'h001c0001);
pulp_write32(axi_m, 32'h44000fa4, 32'h001c0002);
pulp_write32(axi_m, 32'h44000fa8, 32'h001c0003);
pulp_write32(axi_m, 32'h44000fac, 32'h001c0004);
pulp_write32(axi_m, 32'h44000fb0, 32'h001c0005);
pulp_write32(axi_m, 32'h44000fb4, 32'h001c0006);
pulp_write32(axi_m, 32'h44000fb8, 32'h001c0007);
pulp_write32(axi_m, 32'h44000fbc, 32'h001c0008);
pulp_write32(axi_m, 32'h44000fc0, 32'h001c0009);
pulp_write32(axi_m, 32'h44000fc4, 32'h001c000a);
pulp_write32(axi_m, 32'h44000fc8, 32'h001c000b);
pulp_write32(axi_m, 32'h44000fcc, 32'h001c000c);
pulp_write32(axi_m, 32'h44000fd0, 32'h001c000d);
pulp_write32(axi_m, 32'h44000fd4, 32'h001c000e);
pulp_write32(axi_m, 32'h44000fd8, 32'h001c000f);

pulp_write32(axi_m, 32'h44000fdc, 32'd29);
pulp_write32(axi_m, 32'h44000fe0, 32'd2);
pulp_write32(axi_m, 32'h44000fe4, 32'h80001a10);
pulp_write32(axi_m, 32'h44001a10, 32'h80001068);
pulp_write32(axi_m, 32'h44001a14, 32'h80001810);
pulp_write32(axi_m, 32'h44001028, 32'h001d0000);
pulp_write32(axi_m, 32'h4400102c, 32'h001d0001);
pulp_write32(axi_m, 32'h44001030, 32'h001d0002);
pulp_write32(axi_m, 32'h44001034, 32'h001d0003);
pulp_write32(axi_m, 32'h44001038, 32'h001d0004);
pulp_write32(axi_m, 32'h4400103c, 32'h001d0005);
pulp_write32(axi_m, 32'h44001040, 32'h001d0006);
pulp_write32(axi_m, 32'h44001044, 32'h001d0007);
pulp_write32(axi_m, 32'h44001048, 32'h001d0008);
pulp_write32(axi_m, 32'h4400104c, 32'h001d0009);
pulp_write32(axi_m, 32'h44001050, 32'h001d000a);
pulp_write32(axi_m, 32'h44001054, 32'h001d000b);
pulp_write32(axi_m, 32'h44001058, 32'h001d000c);
pulp_write32(axi_m, 32'h4400105c, 32'h001d000d);
pulp_write32(axi_m, 32'h44001060, 32'h001d000e);
pulp_write32(axi_m, 32'h44001064, 32'h001d000f);

pulp_write32(axi_m, 32'h44001068, 32'd30);
pulp_write32(axi_m, 32'h4400106c, 32'd1);
pulp_write32(axi_m, 32'h44001070, 32'h80001a18);
pulp_write32(axi_m, 32'h44001a18, 32'h80001324);
pulp_write32(axi_m, 32'h440010b4, 32'h001e0000);
pulp_write32(axi_m, 32'h440010b8, 32'h001e0001);
pulp_write32(axi_m, 32'h440010bc, 32'h001e0002);
pulp_write32(axi_m, 32'h440010c0, 32'h001e0003);
pulp_write32(axi_m, 32'h440010c4, 32'h001e0004);
pulp_write32(axi_m, 32'h440010c8, 32'h001e0005);
pulp_write32(axi_m, 32'h440010cc, 32'h001e0006);
pulp_write32(axi_m, 32'h440010d0, 32'h001e0007);
pulp_write32(axi_m, 32'h440010d4, 32'h001e0008);
pulp_write32(axi_m, 32'h440010d8, 32'h001e0009);
pulp_write32(axi_m, 32'h440010dc, 32'h001e000a);
pulp_write32(axi_m, 32'h440010e0, 32'h001e000b);
pulp_write32(axi_m, 32'h440010e4, 32'h001e000c);
pulp_write32(axi_m, 32'h440010e8, 32'h001e000d);
pulp_write32(axi_m, 32'h440010ec, 32'h001e000e);
pulp_write32(axi_m, 32'h440010f0, 32'h001e000f);

pulp_write32(axi_m, 32'h440010f4, 32'd31);
pulp_write32(axi_m, 32'h440010f8, 32'd2);
pulp_write32(axi_m, 32'h440010fc, 32'h80001a20);
pulp_write32(axi_m, 32'h44001a20, 32'h80001180);
pulp_write32(axi_m, 32'h44001a24, 32'h80001324);
pulp_write32(axi_m, 32'h44001140, 32'h001f0000);
pulp_write32(axi_m, 32'h44001144, 32'h001f0001);
pulp_write32(axi_m, 32'h44001148, 32'h001f0002);
pulp_write32(axi_m, 32'h4400114c, 32'h001f0003);
pulp_write32(axi_m, 32'h44001150, 32'h001f0004);
pulp_write32(axi_m, 32'h44001154, 32'h001f0005);
pulp_write32(axi_m, 32'h44001158, 32'h001f0006);
pulp_write32(axi_m, 32'h4400115c, 32'h001f0007);
pulp_write32(axi_m, 32'h44001160, 32'h001f0008);
pulp_write32(axi_m, 32'h44001164, 32'h001f0009);
pulp_write32(axi_m, 32'h44001168, 32'h001f000a);
pulp_write32(axi_m, 32'h4400116c, 32'h001f000b);
pulp_write32(axi_m, 32'h44001170, 32'h001f000c);
pulp_write32(axi_m, 32'h44001174, 32'h001f000d);
pulp_write32(axi_m, 32'h44001178, 32'h001f000e);
pulp_write32(axi_m, 32'h4400117c, 32'h001f000f);

pulp_write32(axi_m, 32'h44001180, 32'd32);
pulp_write32(axi_m, 32'h44001184, 32'd2);
pulp_write32(axi_m, 32'h44001188, 32'h80001a28);
pulp_write32(axi_m, 32'h44001a28, 32'h8000120c);
pulp_write32(axi_m, 32'h44001a2c, 32'h800016f8);
pulp_write32(axi_m, 32'h440011cc, 32'h00200000);
pulp_write32(axi_m, 32'h440011d0, 32'h00200001);
pulp_write32(axi_m, 32'h440011d4, 32'h00200002);
pulp_write32(axi_m, 32'h440011d8, 32'h00200003);
pulp_write32(axi_m, 32'h440011dc, 32'h00200004);
pulp_write32(axi_m, 32'h440011e0, 32'h00200005);
pulp_write32(axi_m, 32'h440011e4, 32'h00200006);
pulp_write32(axi_m, 32'h440011e8, 32'h00200007);
pulp_write32(axi_m, 32'h440011ec, 32'h00200008);
pulp_write32(axi_m, 32'h440011f0, 32'h00200009);
pulp_write32(axi_m, 32'h440011f4, 32'h0020000a);
pulp_write32(axi_m, 32'h440011f8, 32'h0020000b);
pulp_write32(axi_m, 32'h440011fc, 32'h0020000c);
pulp_write32(axi_m, 32'h44001200, 32'h0020000d);
pulp_write32(axi_m, 32'h44001204, 32'h0020000e);
pulp_write32(axi_m, 32'h44001208, 32'h0020000f);

pulp_write32(axi_m, 32'h4400120c, 32'd33);
pulp_write32(axi_m, 32'h44001210, 32'd1);
pulp_write32(axi_m, 32'h44001214, 32'h80001a30);
pulp_write32(axi_m, 32'h44001a30, 32'h80001784);
pulp_write32(axi_m, 32'h44001258, 32'h00210000);
pulp_write32(axi_m, 32'h4400125c, 32'h00210001);
pulp_write32(axi_m, 32'h44001260, 32'h00210002);
pulp_write32(axi_m, 32'h44001264, 32'h00210003);
pulp_write32(axi_m, 32'h44001268, 32'h00210004);
pulp_write32(axi_m, 32'h4400126c, 32'h00210005);
pulp_write32(axi_m, 32'h44001270, 32'h00210006);
pulp_write32(axi_m, 32'h44001274, 32'h00210007);
pulp_write32(axi_m, 32'h44001278, 32'h00210008);
pulp_write32(axi_m, 32'h4400127c, 32'h00210009);
pulp_write32(axi_m, 32'h44001280, 32'h0021000a);
pulp_write32(axi_m, 32'h44001284, 32'h0021000b);
pulp_write32(axi_m, 32'h44001288, 32'h0021000c);
pulp_write32(axi_m, 32'h4400128c, 32'h0021000d);
pulp_write32(axi_m, 32'h44001290, 32'h0021000e);
pulp_write32(axi_m, 32'h44001294, 32'h0021000f);

pulp_write32(axi_m, 32'h44001298, 32'd34);
pulp_write32(axi_m, 32'h4400129c, 32'd1);
pulp_write32(axi_m, 32'h440012a0, 32'h80001a38);
pulp_write32(axi_m, 32'h44001a38, 32'h800013b0);
pulp_write32(axi_m, 32'h440012e4, 32'h00220000);
pulp_write32(axi_m, 32'h440012e8, 32'h00220001);
pulp_write32(axi_m, 32'h440012ec, 32'h00220002);
pulp_write32(axi_m, 32'h440012f0, 32'h00220003);
pulp_write32(axi_m, 32'h440012f4, 32'h00220004);
pulp_write32(axi_m, 32'h440012f8, 32'h00220005);
pulp_write32(axi_m, 32'h440012fc, 32'h00220006);
pulp_write32(axi_m, 32'h44001300, 32'h00220007);
pulp_write32(axi_m, 32'h44001304, 32'h00220008);
pulp_write32(axi_m, 32'h44001308, 32'h00220009);
pulp_write32(axi_m, 32'h4400130c, 32'h0022000a);
pulp_write32(axi_m, 32'h44001310, 32'h0022000b);
pulp_write32(axi_m, 32'h44001314, 32'h0022000c);
pulp_write32(axi_m, 32'h44001318, 32'h0022000d);
pulp_write32(axi_m, 32'h4400131c, 32'h0022000e);
pulp_write32(axi_m, 32'h44001320, 32'h0022000f);

pulp_write32(axi_m, 32'h44001324, 32'd35);
pulp_write32(axi_m, 32'h44001328, 32'd1);
pulp_write32(axi_m, 32'h4400132c, 32'h80001a40);
pulp_write32(axi_m, 32'h44001a40, 32'h8000143c);
pulp_write32(axi_m, 32'h44001370, 32'h00230000);
pulp_write32(axi_m, 32'h44001374, 32'h00230001);
pulp_write32(axi_m, 32'h44001378, 32'h00230002);
pulp_write32(axi_m, 32'h4400137c, 32'h00230003);
pulp_write32(axi_m, 32'h44001380, 32'h00230004);
pulp_write32(axi_m, 32'h44001384, 32'h00230005);
pulp_write32(axi_m, 32'h44001388, 32'h00230006);
pulp_write32(axi_m, 32'h4400138c, 32'h00230007);
pulp_write32(axi_m, 32'h44001390, 32'h00230008);
pulp_write32(axi_m, 32'h44001394, 32'h00230009);
pulp_write32(axi_m, 32'h44001398, 32'h0023000a);
pulp_write32(axi_m, 32'h4400139c, 32'h0023000b);
pulp_write32(axi_m, 32'h440013a0, 32'h0023000c);
pulp_write32(axi_m, 32'h440013a4, 32'h0023000d);
pulp_write32(axi_m, 32'h440013a8, 32'h0023000e);
pulp_write32(axi_m, 32'h440013ac, 32'h0023000f);

pulp_write32(axi_m, 32'h440013b0, 32'd36);
pulp_write32(axi_m, 32'h440013b4, 32'd2);
pulp_write32(axi_m, 32'h440013b8, 32'h80001a48);
pulp_write32(axi_m, 32'h44001a48, 32'h800014c8);
pulp_write32(axi_m, 32'h44001a4c, 32'h80001554);
pulp_write32(axi_m, 32'h440013fc, 32'h00240000);
pulp_write32(axi_m, 32'h44001400, 32'h00240001);
pulp_write32(axi_m, 32'h44001404, 32'h00240002);
pulp_write32(axi_m, 32'h44001408, 32'h00240003);
pulp_write32(axi_m, 32'h4400140c, 32'h00240004);
pulp_write32(axi_m, 32'h44001410, 32'h00240005);
pulp_write32(axi_m, 32'h44001414, 32'h00240006);
pulp_write32(axi_m, 32'h44001418, 32'h00240007);
pulp_write32(axi_m, 32'h4400141c, 32'h00240008);
pulp_write32(axi_m, 32'h44001420, 32'h00240009);
pulp_write32(axi_m, 32'h44001424, 32'h0024000a);
pulp_write32(axi_m, 32'h44001428, 32'h0024000b);
pulp_write32(axi_m, 32'h4400142c, 32'h0024000c);
pulp_write32(axi_m, 32'h44001430, 32'h0024000d);
pulp_write32(axi_m, 32'h44001434, 32'h0024000e);
pulp_write32(axi_m, 32'h44001438, 32'h0024000f);

pulp_write32(axi_m, 32'h4400143c, 32'd37);
pulp_write32(axi_m, 32'h44001440, 32'd2);
pulp_write32(axi_m, 32'h44001444, 32'h80001a50);
pulp_write32(axi_m, 32'h44001a50, 32'h800016f8);
pulp_write32(axi_m, 32'h44001a54, 32'h80001810);
pulp_write32(axi_m, 32'h44001488, 32'h00250000);
pulp_write32(axi_m, 32'h4400148c, 32'h00250001);
pulp_write32(axi_m, 32'h44001490, 32'h00250002);
pulp_write32(axi_m, 32'h44001494, 32'h00250003);
pulp_write32(axi_m, 32'h44001498, 32'h00250004);
pulp_write32(axi_m, 32'h4400149c, 32'h00250005);
pulp_write32(axi_m, 32'h440014a0, 32'h00250006);
pulp_write32(axi_m, 32'h440014a4, 32'h00250007);
pulp_write32(axi_m, 32'h440014a8, 32'h00250008);
pulp_write32(axi_m, 32'h440014ac, 32'h00250009);
pulp_write32(axi_m, 32'h440014b0, 32'h0025000a);
pulp_write32(axi_m, 32'h440014b4, 32'h0025000b);
pulp_write32(axi_m, 32'h440014b8, 32'h0025000c);
pulp_write32(axi_m, 32'h440014bc, 32'h0025000d);
pulp_write32(axi_m, 32'h440014c0, 32'h0025000e);
pulp_write32(axi_m, 32'h440014c4, 32'h0025000f);

pulp_write32(axi_m, 32'h440014c8, 32'd38);
pulp_write32(axi_m, 32'h440014cc, 32'd1);
pulp_write32(axi_m, 32'h440014d0, 32'h80001a58);
pulp_write32(axi_m, 32'h44001a58, 32'h800015e0);
pulp_write32(axi_m, 32'h44001514, 32'h00260000);
pulp_write32(axi_m, 32'h44001518, 32'h00260001);
pulp_write32(axi_m, 32'h4400151c, 32'h00260002);
pulp_write32(axi_m, 32'h44001520, 32'h00260003);
pulp_write32(axi_m, 32'h44001524, 32'h00260004);
pulp_write32(axi_m, 32'h44001528, 32'h00260005);
pulp_write32(axi_m, 32'h4400152c, 32'h00260006);
pulp_write32(axi_m, 32'h44001530, 32'h00260007);
pulp_write32(axi_m, 32'h44001534, 32'h00260008);
pulp_write32(axi_m, 32'h44001538, 32'h00260009);
pulp_write32(axi_m, 32'h4400153c, 32'h0026000a);
pulp_write32(axi_m, 32'h44001540, 32'h0026000b);
pulp_write32(axi_m, 32'h44001544, 32'h0026000c);
pulp_write32(axi_m, 32'h44001548, 32'h0026000d);
pulp_write32(axi_m, 32'h4400154c, 32'h0026000e);
pulp_write32(axi_m, 32'h44001550, 32'h0026000f);

pulp_write32(axi_m, 32'h44001554, 32'd39);
pulp_write32(axi_m, 32'h44001558, 32'd1);
pulp_write32(axi_m, 32'h4400155c, 32'h80001a60);
pulp_write32(axi_m, 32'h44001a60, 32'h8000166c);
pulp_write32(axi_m, 32'h440015a0, 32'h00270000);
pulp_write32(axi_m, 32'h440015a4, 32'h00270001);
pulp_write32(axi_m, 32'h440015a8, 32'h00270002);
pulp_write32(axi_m, 32'h440015ac, 32'h00270003);
pulp_write32(axi_m, 32'h440015b0, 32'h00270004);
pulp_write32(axi_m, 32'h440015b4, 32'h00270005);
pulp_write32(axi_m, 32'h440015b8, 32'h00270006);
pulp_write32(axi_m, 32'h440015bc, 32'h00270007);
pulp_write32(axi_m, 32'h440015c0, 32'h00270008);
pulp_write32(axi_m, 32'h440015c4, 32'h00270009);
pulp_write32(axi_m, 32'h440015c8, 32'h0027000a);
pulp_write32(axi_m, 32'h440015cc, 32'h0027000b);
pulp_write32(axi_m, 32'h440015d0, 32'h0027000c);
pulp_write32(axi_m, 32'h440015d4, 32'h0027000d);
pulp_write32(axi_m, 32'h440015d8, 32'h0027000e);
pulp_write32(axi_m, 32'h440015dc, 32'h0027000f);

pulp_write32(axi_m, 32'h440015e0, 32'd40);
pulp_write32(axi_m, 32'h440015e4, 32'd1);
pulp_write32(axi_m, 32'h440015e8, 32'h80001a68);
pulp_write32(axi_m, 32'h44001a68, 32'h8000166c);
pulp_write32(axi_m, 32'h4400162c, 32'h00280000);
pulp_write32(axi_m, 32'h44001630, 32'h00280001);
pulp_write32(axi_m, 32'h44001634, 32'h00280002);
pulp_write32(axi_m, 32'h44001638, 32'h00280003);
pulp_write32(axi_m, 32'h4400163c, 32'h00280004);
pulp_write32(axi_m, 32'h44001640, 32'h00280005);
pulp_write32(axi_m, 32'h44001644, 32'h00280006);
pulp_write32(axi_m, 32'h44001648, 32'h00280007);
pulp_write32(axi_m, 32'h4400164c, 32'h00280008);
pulp_write32(axi_m, 32'h44001650, 32'h00280009);
pulp_write32(axi_m, 32'h44001654, 32'h0028000a);
pulp_write32(axi_m, 32'h44001658, 32'h0028000b);
pulp_write32(axi_m, 32'h4400165c, 32'h0028000c);
pulp_write32(axi_m, 32'h44001660, 32'h0028000d);
pulp_write32(axi_m, 32'h44001664, 32'h0028000e);
pulp_write32(axi_m, 32'h44001668, 32'h0028000f);

pulp_write32(axi_m, 32'h4400166c, 32'd41);
pulp_write32(axi_m, 32'h44001670, 32'd0);
pulp_write32(axi_m, 32'h440016b8, 32'h00290000);
pulp_write32(axi_m, 32'h440016bc, 32'h00290001);
pulp_write32(axi_m, 32'h440016c0, 32'h00290002);
pulp_write32(axi_m, 32'h440016c4, 32'h00290003);
pulp_write32(axi_m, 32'h440016c8, 32'h00290004);
pulp_write32(axi_m, 32'h440016cc, 32'h00290005);
pulp_write32(axi_m, 32'h440016d0, 32'h00290006);
pulp_write32(axi_m, 32'h440016d4, 32'h00290007);
pulp_write32(axi_m, 32'h440016d8, 32'h00290008);
pulp_write32(axi_m, 32'h440016dc, 32'h00290009);
pulp_write32(axi_m, 32'h440016e0, 32'h0029000a);
pulp_write32(axi_m, 32'h440016e4, 32'h0029000b);
pulp_write32(axi_m, 32'h440016e8, 32'h0029000c);
pulp_write32(axi_m, 32'h440016ec, 32'h0029000d);
pulp_write32(axi_m, 32'h440016f0, 32'h0029000e);
pulp_write32(axi_m, 32'h440016f4, 32'h0029000f);

pulp_write32(axi_m, 32'h440016f8, 32'd42);
pulp_write32(axi_m, 32'h440016fc, 32'd1);
pulp_write32(axi_m, 32'h44001700, 32'h80001a70);
pulp_write32(axi_m, 32'h44001a70, 32'h80001784);
pulp_write32(axi_m, 32'h44001744, 32'h002a0000);
pulp_write32(axi_m, 32'h44001748, 32'h002a0001);
pulp_write32(axi_m, 32'h4400174c, 32'h002a0002);
pulp_write32(axi_m, 32'h44001750, 32'h002a0003);
pulp_write32(axi_m, 32'h44001754, 32'h002a0004);
pulp_write32(axi_m, 32'h44001758, 32'h002a0005);
pulp_write32(axi_m, 32'h4400175c, 32'h002a0006);
pulp_write32(axi_m, 32'h44001760, 32'h002a0007);
pulp_write32(axi_m, 32'h44001764, 32'h002a0008);
pulp_write32(axi_m, 32'h44001768, 32'h002a0009);
pulp_write32(axi_m, 32'h4400176c, 32'h002a000a);
pulp_write32(axi_m, 32'h44001770, 32'h002a000b);
pulp_write32(axi_m, 32'h44001774, 32'h002a000c);
pulp_write32(axi_m, 32'h44001778, 32'h002a000d);
pulp_write32(axi_m, 32'h4400177c, 32'h002a000e);
pulp_write32(axi_m, 32'h44001780, 32'h002a000f);

pulp_write32(axi_m, 32'h44001784, 32'd43);
pulp_write32(axi_m, 32'h44001788, 32'd1);
pulp_write32(axi_m, 32'h4400178c, 32'h80001a78);
pulp_write32(axi_m, 32'h44001a78, 32'h8000189c);
pulp_write32(axi_m, 32'h440017d0, 32'h002b0000);
pulp_write32(axi_m, 32'h440017d4, 32'h002b0001);
pulp_write32(axi_m, 32'h440017d8, 32'h002b0002);
pulp_write32(axi_m, 32'h440017dc, 32'h002b0003);
pulp_write32(axi_m, 32'h440017e0, 32'h002b0004);
pulp_write32(axi_m, 32'h440017e4, 32'h002b0005);
pulp_write32(axi_m, 32'h440017e8, 32'h002b0006);
pulp_write32(axi_m, 32'h440017ec, 32'h002b0007);
pulp_write32(axi_m, 32'h440017f0, 32'h002b0008);
pulp_write32(axi_m, 32'h440017f4, 32'h002b0009);
pulp_write32(axi_m, 32'h440017f8, 32'h002b000a);
pulp_write32(axi_m, 32'h440017fc, 32'h002b000b);
pulp_write32(axi_m, 32'h44001800, 32'h002b000c);
pulp_write32(axi_m, 32'h44001804, 32'h002b000d);
pulp_write32(axi_m, 32'h44001808, 32'h002b000e);
pulp_write32(axi_m, 32'h4400180c, 32'h002b000f);

pulp_write32(axi_m, 32'h44001810, 32'd44);
pulp_write32(axi_m, 32'h44001814, 32'd1);
pulp_write32(axi_m, 32'h44001818, 32'h80001a80);
pulp_write32(axi_m, 32'h44001a80, 32'h8000189c);
pulp_write32(axi_m, 32'h4400185c, 32'h002c0000);
pulp_write32(axi_m, 32'h44001860, 32'h002c0001);
pulp_write32(axi_m, 32'h44001864, 32'h002c0002);
pulp_write32(axi_m, 32'h44001868, 32'h002c0003);
pulp_write32(axi_m, 32'h4400186c, 32'h002c0004);
pulp_write32(axi_m, 32'h44001870, 32'h002c0005);
pulp_write32(axi_m, 32'h44001874, 32'h002c0006);
pulp_write32(axi_m, 32'h44001878, 32'h002c0007);
pulp_write32(axi_m, 32'h4400187c, 32'h002c0008);
pulp_write32(axi_m, 32'h44001880, 32'h002c0009);
pulp_write32(axi_m, 32'h44001884, 32'h002c000a);
pulp_write32(axi_m, 32'h44001888, 32'h002c000b);
pulp_write32(axi_m, 32'h4400188c, 32'h002c000c);
pulp_write32(axi_m, 32'h44001890, 32'h002c000d);
pulp_write32(axi_m, 32'h44001894, 32'h002c000e);
pulp_write32(axi_m, 32'h44001898, 32'h002c000f);

pulp_write32(axi_m, 32'h4400189c, 32'd45);
pulp_write32(axi_m, 32'h440018a0, 32'd0);
pulp_write32(axi_m, 32'h440018e8, 32'h002d0000);
pulp_write32(axi_m, 32'h440018ec, 32'h002d0001);
pulp_write32(axi_m, 32'h440018f0, 32'h002d0002);
pulp_write32(axi_m, 32'h440018f4, 32'h002d0003);
pulp_write32(axi_m, 32'h440018f8, 32'h002d0004);
pulp_write32(axi_m, 32'h440018fc, 32'h002d0005);
pulp_write32(axi_m, 32'h44001900, 32'h002d0006);
pulp_write32(axi_m, 32'h44001904, 32'h002d0007);
pulp_write32(axi_m, 32'h44001908, 32'h002d0008);
pulp_write32(axi_m, 32'h4400190c, 32'h002d0009);
pulp_write32(axi_m, 32'h44001910, 32'h002d000a);
pulp_write32(axi_m, 32'h44001914, 32'h002d000b);
pulp_write32(axi_m, 32'h44001918, 32'h002d000c);
pulp_write32(axi_m, 32'h4400191c, 32'h002d000d);
pulp_write32(axi_m, 32'h44001920, 32'h002d000e);
pulp_write32(axi_m, 32'h44001924, 32'h002d000f);

