pulp_write32(axi_m, 32'ha4000000, 32'd0);
pulp_write32(axi_m, 32'ha4000004, 32'd3);
pulp_write32(axi_m, 32'ha4000008, 32'h80001928);
pulp_write32(axi_m, 32'ha4001928, 32'h80000578);
pulp_write32(axi_m, 32'ha400192c, 32'h80000604);
pulp_write32(axi_m, 32'ha4001930, 32'h80000690);
pulp_write32(axi_m, 32'ha400004c, 32'h00000000);
pulp_write32(axi_m, 32'ha4000050, 32'h00000001);
pulp_write32(axi_m, 32'ha4000054, 32'h00000002);
pulp_write32(axi_m, 32'ha4000058, 32'h00000003);
pulp_write32(axi_m, 32'ha400005c, 32'h00000004);
pulp_write32(axi_m, 32'ha4000060, 32'h00000005);
pulp_write32(axi_m, 32'ha4000064, 32'h00000006);
pulp_write32(axi_m, 32'ha4000068, 32'h00000007);
pulp_write32(axi_m, 32'ha400006c, 32'h00000008);
pulp_write32(axi_m, 32'ha4000070, 32'h00000009);
pulp_write32(axi_m, 32'ha4000074, 32'h0000000a);
pulp_write32(axi_m, 32'ha4000078, 32'h0000000b);
pulp_write32(axi_m, 32'ha400007c, 32'h0000000c);
pulp_write32(axi_m, 32'ha4000080, 32'h0000000d);
pulp_write32(axi_m, 32'ha4000084, 32'h0000000e);
pulp_write32(axi_m, 32'ha4000088, 32'h0000000f);

pulp_write32(axi_m, 32'ha400008c, 32'd1);
pulp_write32(axi_m, 32'ha4000090, 32'd3);
pulp_write32(axi_m, 32'ha4000094, 32'h80001938);
pulp_write32(axi_m, 32'ha4001938, 32'h80000118);
pulp_write32(axi_m, 32'ha400193c, 32'h800003d4);
pulp_write32(axi_m, 32'ha4001940, 32'h80000a64);
pulp_write32(axi_m, 32'ha40000d8, 32'h00010000);
pulp_write32(axi_m, 32'ha40000dc, 32'h00010001);
pulp_write32(axi_m, 32'ha40000e0, 32'h00010002);
pulp_write32(axi_m, 32'ha40000e4, 32'h00010003);
pulp_write32(axi_m, 32'ha40000e8, 32'h00010004);
pulp_write32(axi_m, 32'ha40000ec, 32'h00010005);
pulp_write32(axi_m, 32'ha40000f0, 32'h00010006);
pulp_write32(axi_m, 32'ha40000f4, 32'h00010007);
pulp_write32(axi_m, 32'ha40000f8, 32'h00010008);
pulp_write32(axi_m, 32'ha40000fc, 32'h00010009);
pulp_write32(axi_m, 32'ha4000100, 32'h0001000a);
pulp_write32(axi_m, 32'ha4000104, 32'h0001000b);
pulp_write32(axi_m, 32'ha4000108, 32'h0001000c);
pulp_write32(axi_m, 32'ha400010c, 32'h0001000d);
pulp_write32(axi_m, 32'ha4000110, 32'h0001000e);
pulp_write32(axi_m, 32'ha4000114, 32'h0001000f);

pulp_write32(axi_m, 32'ha4000118, 32'd2);
pulp_write32(axi_m, 32'ha400011c, 32'd2);
pulp_write32(axi_m, 32'ha4000120, 32'h80001948);
pulp_write32(axi_m, 32'ha4001948, 32'h800001a4);
pulp_write32(axi_m, 32'ha400194c, 32'h8000166c);
pulp_write32(axi_m, 32'ha4000164, 32'h00020000);
pulp_write32(axi_m, 32'ha4000168, 32'h00020001);
pulp_write32(axi_m, 32'ha400016c, 32'h00020002);
pulp_write32(axi_m, 32'ha4000170, 32'h00020003);
pulp_write32(axi_m, 32'ha4000174, 32'h00020004);
pulp_write32(axi_m, 32'ha4000178, 32'h00020005);
pulp_write32(axi_m, 32'ha400017c, 32'h00020006);
pulp_write32(axi_m, 32'ha4000180, 32'h00020007);
pulp_write32(axi_m, 32'ha4000184, 32'h00020008);
pulp_write32(axi_m, 32'ha4000188, 32'h00020009);
pulp_write32(axi_m, 32'ha400018c, 32'h0002000a);
pulp_write32(axi_m, 32'ha4000190, 32'h0002000b);
pulp_write32(axi_m, 32'ha4000194, 32'h0002000c);
pulp_write32(axi_m, 32'ha4000198, 32'h0002000d);
pulp_write32(axi_m, 32'ha400019c, 32'h0002000e);
pulp_write32(axi_m, 32'ha40001a0, 32'h0002000f);

pulp_write32(axi_m, 32'ha40001a4, 32'd3);
pulp_write32(axi_m, 32'ha40001a8, 32'd2);
pulp_write32(axi_m, 32'ha40001ac, 32'h80001950);
pulp_write32(axi_m, 32'ha4001950, 32'h80000230);
pulp_write32(axi_m, 32'ha4001954, 32'h80000ec4);
pulp_write32(axi_m, 32'ha40001f0, 32'h00030000);
pulp_write32(axi_m, 32'ha40001f4, 32'h00030001);
pulp_write32(axi_m, 32'ha40001f8, 32'h00030002);
pulp_write32(axi_m, 32'ha40001fc, 32'h00030003);
pulp_write32(axi_m, 32'ha4000200, 32'h00030004);
pulp_write32(axi_m, 32'ha4000204, 32'h00030005);
pulp_write32(axi_m, 32'ha4000208, 32'h00030006);
pulp_write32(axi_m, 32'ha400020c, 32'h00030007);
pulp_write32(axi_m, 32'ha4000210, 32'h00030008);
pulp_write32(axi_m, 32'ha4000214, 32'h00030009);
pulp_write32(axi_m, 32'ha4000218, 32'h0003000a);
pulp_write32(axi_m, 32'ha400021c, 32'h0003000b);
pulp_write32(axi_m, 32'ha4000220, 32'h0003000c);
pulp_write32(axi_m, 32'ha4000224, 32'h0003000d);
pulp_write32(axi_m, 32'ha4000228, 32'h0003000e);
pulp_write32(axi_m, 32'ha400022c, 32'h0003000f);

pulp_write32(axi_m, 32'ha4000230, 32'd4);
pulp_write32(axi_m, 32'ha4000234, 32'd2);
pulp_write32(axi_m, 32'ha4000238, 32'h80001958);
pulp_write32(axi_m, 32'ha4001958, 32'h800002bc);
pulp_write32(axi_m, 32'ha400195c, 32'h8000120c);
pulp_write32(axi_m, 32'ha400027c, 32'h00040000);
pulp_write32(axi_m, 32'ha4000280, 32'h00040001);
pulp_write32(axi_m, 32'ha4000284, 32'h00040002);
pulp_write32(axi_m, 32'ha4000288, 32'h00040003);
pulp_write32(axi_m, 32'ha400028c, 32'h00040004);
pulp_write32(axi_m, 32'ha4000290, 32'h00040005);
pulp_write32(axi_m, 32'ha4000294, 32'h00040006);
pulp_write32(axi_m, 32'ha4000298, 32'h00040007);
pulp_write32(axi_m, 32'ha400029c, 32'h00040008);
pulp_write32(axi_m, 32'ha40002a0, 32'h00040009);
pulp_write32(axi_m, 32'ha40002a4, 32'h0004000a);
pulp_write32(axi_m, 32'ha40002a8, 32'h0004000b);
pulp_write32(axi_m, 32'ha40002ac, 32'h0004000c);
pulp_write32(axi_m, 32'ha40002b0, 32'h0004000d);
pulp_write32(axi_m, 32'ha40002b4, 32'h0004000e);
pulp_write32(axi_m, 32'ha40002b8, 32'h0004000f);

pulp_write32(axi_m, 32'ha40002bc, 32'd5);
pulp_write32(axi_m, 32'ha40002c0, 32'd2);
pulp_write32(axi_m, 32'ha40002c4, 32'h80001960);
pulp_write32(axi_m, 32'ha4001960, 32'h80000348);
pulp_write32(axi_m, 32'ha4001964, 32'h8000189c);
pulp_write32(axi_m, 32'ha4000308, 32'h00050000);
pulp_write32(axi_m, 32'ha400030c, 32'h00050001);
pulp_write32(axi_m, 32'ha4000310, 32'h00050002);
pulp_write32(axi_m, 32'ha4000314, 32'h00050003);
pulp_write32(axi_m, 32'ha4000318, 32'h00050004);
pulp_write32(axi_m, 32'ha400031c, 32'h00050005);
pulp_write32(axi_m, 32'ha4000320, 32'h00050006);
pulp_write32(axi_m, 32'ha4000324, 32'h00050007);
pulp_write32(axi_m, 32'ha4000328, 32'h00050008);
pulp_write32(axi_m, 32'ha400032c, 32'h00050009);
pulp_write32(axi_m, 32'ha4000330, 32'h0005000a);
pulp_write32(axi_m, 32'ha4000334, 32'h0005000b);
pulp_write32(axi_m, 32'ha4000338, 32'h0005000c);
pulp_write32(axi_m, 32'ha400033c, 32'h0005000d);
pulp_write32(axi_m, 32'ha4000340, 32'h0005000e);
pulp_write32(axi_m, 32'ha4000344, 32'h0005000f);

pulp_write32(axi_m, 32'ha4000348, 32'd6);
pulp_write32(axi_m, 32'ha400034c, 32'd2);
pulp_write32(axi_m, 32'ha4000350, 32'h80001968);
pulp_write32(axi_m, 32'ha4001968, 32'h800004ec);
pulp_write32(axi_m, 32'ha400196c, 32'h80000fdc);
pulp_write32(axi_m, 32'ha4000394, 32'h00060000);
pulp_write32(axi_m, 32'ha4000398, 32'h00060001);
pulp_write32(axi_m, 32'ha400039c, 32'h00060002);
pulp_write32(axi_m, 32'ha40003a0, 32'h00060003);
pulp_write32(axi_m, 32'ha40003a4, 32'h00060004);
pulp_write32(axi_m, 32'ha40003a8, 32'h00060005);
pulp_write32(axi_m, 32'ha40003ac, 32'h00060006);
pulp_write32(axi_m, 32'ha40003b0, 32'h00060007);
pulp_write32(axi_m, 32'ha40003b4, 32'h00060008);
pulp_write32(axi_m, 32'ha40003b8, 32'h00060009);
pulp_write32(axi_m, 32'ha40003bc, 32'h0006000a);
pulp_write32(axi_m, 32'ha40003c0, 32'h0006000b);
pulp_write32(axi_m, 32'ha40003c4, 32'h0006000c);
pulp_write32(axi_m, 32'ha40003c8, 32'h0006000d);
pulp_write32(axi_m, 32'ha40003cc, 32'h0006000e);
pulp_write32(axi_m, 32'ha40003d0, 32'h0006000f);

pulp_write32(axi_m, 32'ha40003d4, 32'd7);
pulp_write32(axi_m, 32'ha40003d8, 32'd2);
pulp_write32(axi_m, 32'ha40003dc, 32'h80001970);
pulp_write32(axi_m, 32'ha4001970, 32'h80000460);
pulp_write32(axi_m, 32'ha4001974, 32'h80000b7c);
pulp_write32(axi_m, 32'ha4000420, 32'h00070000);
pulp_write32(axi_m, 32'ha4000424, 32'h00070001);
pulp_write32(axi_m, 32'ha4000428, 32'h00070002);
pulp_write32(axi_m, 32'ha400042c, 32'h00070003);
pulp_write32(axi_m, 32'ha4000430, 32'h00070004);
pulp_write32(axi_m, 32'ha4000434, 32'h00070005);
pulp_write32(axi_m, 32'ha4000438, 32'h00070006);
pulp_write32(axi_m, 32'ha400043c, 32'h00070007);
pulp_write32(axi_m, 32'ha4000440, 32'h00070008);
pulp_write32(axi_m, 32'ha4000444, 32'h00070009);
pulp_write32(axi_m, 32'ha4000448, 32'h0007000a);
pulp_write32(axi_m, 32'ha400044c, 32'h0007000b);
pulp_write32(axi_m, 32'ha4000450, 32'h0007000c);
pulp_write32(axi_m, 32'ha4000454, 32'h0007000d);
pulp_write32(axi_m, 32'ha4000458, 32'h0007000e);
pulp_write32(axi_m, 32'ha400045c, 32'h0007000f);

pulp_write32(axi_m, 32'ha4000460, 32'd8);
pulp_write32(axi_m, 32'ha4000464, 32'd2);
pulp_write32(axi_m, 32'ha4000468, 32'h80001978);
pulp_write32(axi_m, 32'ha4001978, 32'h800004ec);
pulp_write32(axi_m, 32'ha400197c, 32'h80000c08);
pulp_write32(axi_m, 32'ha40004ac, 32'h00080000);
pulp_write32(axi_m, 32'ha40004b0, 32'h00080001);
pulp_write32(axi_m, 32'ha40004b4, 32'h00080002);
pulp_write32(axi_m, 32'ha40004b8, 32'h00080003);
pulp_write32(axi_m, 32'ha40004bc, 32'h00080004);
pulp_write32(axi_m, 32'ha40004c0, 32'h00080005);
pulp_write32(axi_m, 32'ha40004c4, 32'h00080006);
pulp_write32(axi_m, 32'ha40004c8, 32'h00080007);
pulp_write32(axi_m, 32'ha40004cc, 32'h00080008);
pulp_write32(axi_m, 32'ha40004d0, 32'h00080009);
pulp_write32(axi_m, 32'ha40004d4, 32'h0008000a);
pulp_write32(axi_m, 32'ha40004d8, 32'h0008000b);
pulp_write32(axi_m, 32'ha40004dc, 32'h0008000c);
pulp_write32(axi_m, 32'ha40004e0, 32'h0008000d);
pulp_write32(axi_m, 32'ha40004e4, 32'h0008000e);
pulp_write32(axi_m, 32'ha40004e8, 32'h0008000f);

pulp_write32(axi_m, 32'ha40004ec, 32'd9);
pulp_write32(axi_m, 32'ha40004f0, 32'd1);
pulp_write32(axi_m, 32'ha40004f4, 32'h80001980);
pulp_write32(axi_m, 32'ha4001980, 32'h80000d20);
pulp_write32(axi_m, 32'ha4000538, 32'h00090000);
pulp_write32(axi_m, 32'ha400053c, 32'h00090001);
pulp_write32(axi_m, 32'ha4000540, 32'h00090002);
pulp_write32(axi_m, 32'ha4000544, 32'h00090003);
pulp_write32(axi_m, 32'ha4000548, 32'h00090004);
pulp_write32(axi_m, 32'ha400054c, 32'h00090005);
pulp_write32(axi_m, 32'ha4000550, 32'h00090006);
pulp_write32(axi_m, 32'ha4000554, 32'h00090007);
pulp_write32(axi_m, 32'ha4000558, 32'h00090008);
pulp_write32(axi_m, 32'ha400055c, 32'h00090009);
pulp_write32(axi_m, 32'ha4000560, 32'h0009000a);
pulp_write32(axi_m, 32'ha4000564, 32'h0009000b);
pulp_write32(axi_m, 32'ha4000568, 32'h0009000c);
pulp_write32(axi_m, 32'ha400056c, 32'h0009000d);
pulp_write32(axi_m, 32'ha4000570, 32'h0009000e);
pulp_write32(axi_m, 32'ha4000574, 32'h0009000f);

pulp_write32(axi_m, 32'ha4000578, 32'd10);
pulp_write32(axi_m, 32'ha400057c, 32'd2);
pulp_write32(axi_m, 32'ha4000580, 32'h80001988);
pulp_write32(axi_m, 32'ha4001988, 32'h8000071c);
pulp_write32(axi_m, 32'ha400198c, 32'h800007a8);
pulp_write32(axi_m, 32'ha40005c4, 32'h000a0000);
pulp_write32(axi_m, 32'ha40005c8, 32'h000a0001);
pulp_write32(axi_m, 32'ha40005cc, 32'h000a0002);
pulp_write32(axi_m, 32'ha40005d0, 32'h000a0003);
pulp_write32(axi_m, 32'ha40005d4, 32'h000a0004);
pulp_write32(axi_m, 32'ha40005d8, 32'h000a0005);
pulp_write32(axi_m, 32'ha40005dc, 32'h000a0006);
pulp_write32(axi_m, 32'ha40005e0, 32'h000a0007);
pulp_write32(axi_m, 32'ha40005e4, 32'h000a0008);
pulp_write32(axi_m, 32'ha40005e8, 32'h000a0009);
pulp_write32(axi_m, 32'ha40005ec, 32'h000a000a);
pulp_write32(axi_m, 32'ha40005f0, 32'h000a000b);
pulp_write32(axi_m, 32'ha40005f4, 32'h000a000c);
pulp_write32(axi_m, 32'ha40005f8, 32'h000a000d);
pulp_write32(axi_m, 32'ha40005fc, 32'h000a000e);
pulp_write32(axi_m, 32'ha4000600, 32'h000a000f);

pulp_write32(axi_m, 32'ha4000604, 32'd11);
pulp_write32(axi_m, 32'ha4000608, 32'd2);
pulp_write32(axi_m, 32'ha400060c, 32'h80001990);
pulp_write32(axi_m, 32'ha4001990, 32'h80000e38);
pulp_write32(axi_m, 32'ha4001994, 32'h80000f50);
pulp_write32(axi_m, 32'ha4000650, 32'h000b0000);
pulp_write32(axi_m, 32'ha4000654, 32'h000b0001);
pulp_write32(axi_m, 32'ha4000658, 32'h000b0002);
pulp_write32(axi_m, 32'ha400065c, 32'h000b0003);
pulp_write32(axi_m, 32'ha4000660, 32'h000b0004);
pulp_write32(axi_m, 32'ha4000664, 32'h000b0005);
pulp_write32(axi_m, 32'ha4000668, 32'h000b0006);
pulp_write32(axi_m, 32'ha400066c, 32'h000b0007);
pulp_write32(axi_m, 32'ha4000670, 32'h000b0008);
pulp_write32(axi_m, 32'ha4000674, 32'h000b0009);
pulp_write32(axi_m, 32'ha4000678, 32'h000b000a);
pulp_write32(axi_m, 32'ha400067c, 32'h000b000b);
pulp_write32(axi_m, 32'ha4000680, 32'h000b000c);
pulp_write32(axi_m, 32'ha4000684, 32'h000b000d);
pulp_write32(axi_m, 32'ha4000688, 32'h000b000e);
pulp_write32(axi_m, 32'ha400068c, 32'h000b000f);

pulp_write32(axi_m, 32'ha4000690, 32'd12);
pulp_write32(axi_m, 32'ha4000694, 32'd2);
pulp_write32(axi_m, 32'ha4000698, 32'h80001998);
pulp_write32(axi_m, 32'ha4001998, 32'h80001068);
pulp_write32(axi_m, 32'ha400199c, 32'h800010f4);
pulp_write32(axi_m, 32'ha40006dc, 32'h000c0000);
pulp_write32(axi_m, 32'ha40006e0, 32'h000c0001);
pulp_write32(axi_m, 32'ha40006e4, 32'h000c0002);
pulp_write32(axi_m, 32'ha40006e8, 32'h000c0003);
pulp_write32(axi_m, 32'ha40006ec, 32'h000c0004);
pulp_write32(axi_m, 32'ha40006f0, 32'h000c0005);
pulp_write32(axi_m, 32'ha40006f4, 32'h000c0006);
pulp_write32(axi_m, 32'ha40006f8, 32'h000c0007);
pulp_write32(axi_m, 32'ha40006fc, 32'h000c0008);
pulp_write32(axi_m, 32'ha4000700, 32'h000c0009);
pulp_write32(axi_m, 32'ha4000704, 32'h000c000a);
pulp_write32(axi_m, 32'ha4000708, 32'h000c000b);
pulp_write32(axi_m, 32'ha400070c, 32'h000c000c);
pulp_write32(axi_m, 32'ha4000710, 32'h000c000d);
pulp_write32(axi_m, 32'ha4000714, 32'h000c000e);
pulp_write32(axi_m, 32'ha4000718, 32'h000c000f);

pulp_write32(axi_m, 32'ha400071c, 32'd13);
pulp_write32(axi_m, 32'ha4000720, 32'd2);
pulp_write32(axi_m, 32'ha4000724, 32'h800019a0);
pulp_write32(axi_m, 32'ha40019a0, 32'h80000834);
pulp_write32(axi_m, 32'ha40019a4, 32'h80000b7c);
pulp_write32(axi_m, 32'ha4000768, 32'h000d0000);
pulp_write32(axi_m, 32'ha400076c, 32'h000d0001);
pulp_write32(axi_m, 32'ha4000770, 32'h000d0002);
pulp_write32(axi_m, 32'ha4000774, 32'h000d0003);
pulp_write32(axi_m, 32'ha4000778, 32'h000d0004);
pulp_write32(axi_m, 32'ha400077c, 32'h000d0005);
pulp_write32(axi_m, 32'ha4000780, 32'h000d0006);
pulp_write32(axi_m, 32'ha4000784, 32'h000d0007);
pulp_write32(axi_m, 32'ha4000788, 32'h000d0008);
pulp_write32(axi_m, 32'ha400078c, 32'h000d0009);
pulp_write32(axi_m, 32'ha4000790, 32'h000d000a);
pulp_write32(axi_m, 32'ha4000794, 32'h000d000b);
pulp_write32(axi_m, 32'ha4000798, 32'h000d000c);
pulp_write32(axi_m, 32'ha400079c, 32'h000d000d);
pulp_write32(axi_m, 32'ha40007a0, 32'h000d000e);
pulp_write32(axi_m, 32'ha40007a4, 32'h000d000f);

pulp_write32(axi_m, 32'ha40007a8, 32'd14);
pulp_write32(axi_m, 32'ha40007ac, 32'd2);
pulp_write32(axi_m, 32'ha40007b0, 32'h800019a8);
pulp_write32(axi_m, 32'ha40019a8, 32'h80000834);
pulp_write32(axi_m, 32'ha40019ac, 32'h800009d8);
pulp_write32(axi_m, 32'ha40007f4, 32'h000e0000);
pulp_write32(axi_m, 32'ha40007f8, 32'h000e0001);
pulp_write32(axi_m, 32'ha40007fc, 32'h000e0002);
pulp_write32(axi_m, 32'ha4000800, 32'h000e0003);
pulp_write32(axi_m, 32'ha4000804, 32'h000e0004);
pulp_write32(axi_m, 32'ha4000808, 32'h000e0005);
pulp_write32(axi_m, 32'ha400080c, 32'h000e0006);
pulp_write32(axi_m, 32'ha4000810, 32'h000e0007);
pulp_write32(axi_m, 32'ha4000814, 32'h000e0008);
pulp_write32(axi_m, 32'ha4000818, 32'h000e0009);
pulp_write32(axi_m, 32'ha400081c, 32'h000e000a);
pulp_write32(axi_m, 32'ha4000820, 32'h000e000b);
pulp_write32(axi_m, 32'ha4000824, 32'h000e000c);
pulp_write32(axi_m, 32'ha4000828, 32'h000e000d);
pulp_write32(axi_m, 32'ha400082c, 32'h000e000e);
pulp_write32(axi_m, 32'ha4000830, 32'h000e000f);

pulp_write32(axi_m, 32'ha4000834, 32'd15);
pulp_write32(axi_m, 32'ha4000838, 32'd1);
pulp_write32(axi_m, 32'ha400083c, 32'h800019b0);
pulp_write32(axi_m, 32'ha40019b0, 32'h800008c0);
pulp_write32(axi_m, 32'ha4000880, 32'h000f0000);
pulp_write32(axi_m, 32'ha4000884, 32'h000f0001);
pulp_write32(axi_m, 32'ha4000888, 32'h000f0002);
pulp_write32(axi_m, 32'ha400088c, 32'h000f0003);
pulp_write32(axi_m, 32'ha4000890, 32'h000f0004);
pulp_write32(axi_m, 32'ha4000894, 32'h000f0005);
pulp_write32(axi_m, 32'ha4000898, 32'h000f0006);
pulp_write32(axi_m, 32'ha400089c, 32'h000f0007);
pulp_write32(axi_m, 32'ha40008a0, 32'h000f0008);
pulp_write32(axi_m, 32'ha40008a4, 32'h000f0009);
pulp_write32(axi_m, 32'ha40008a8, 32'h000f000a);
pulp_write32(axi_m, 32'ha40008ac, 32'h000f000b);
pulp_write32(axi_m, 32'ha40008b0, 32'h000f000c);
pulp_write32(axi_m, 32'ha40008b4, 32'h000f000d);
pulp_write32(axi_m, 32'ha40008b8, 32'h000f000e);
pulp_write32(axi_m, 32'ha40008bc, 32'h000f000f);

pulp_write32(axi_m, 32'ha40008c0, 32'd16);
pulp_write32(axi_m, 32'ha40008c4, 32'd2);
pulp_write32(axi_m, 32'ha40008c8, 32'h800019b8);
pulp_write32(axi_m, 32'ha40019b8, 32'h8000094c);
pulp_write32(axi_m, 32'ha40019bc, 32'h80000af0);
pulp_write32(axi_m, 32'ha400090c, 32'h00100000);
pulp_write32(axi_m, 32'ha4000910, 32'h00100001);
pulp_write32(axi_m, 32'ha4000914, 32'h00100002);
pulp_write32(axi_m, 32'ha4000918, 32'h00100003);
pulp_write32(axi_m, 32'ha400091c, 32'h00100004);
pulp_write32(axi_m, 32'ha4000920, 32'h00100005);
pulp_write32(axi_m, 32'ha4000924, 32'h00100006);
pulp_write32(axi_m, 32'ha4000928, 32'h00100007);
pulp_write32(axi_m, 32'ha400092c, 32'h00100008);
pulp_write32(axi_m, 32'ha4000930, 32'h00100009);
pulp_write32(axi_m, 32'ha4000934, 32'h0010000a);
pulp_write32(axi_m, 32'ha4000938, 32'h0010000b);
pulp_write32(axi_m, 32'ha400093c, 32'h0010000c);
pulp_write32(axi_m, 32'ha4000940, 32'h0010000d);
pulp_write32(axi_m, 32'ha4000944, 32'h0010000e);
pulp_write32(axi_m, 32'ha4000948, 32'h0010000f);

pulp_write32(axi_m, 32'ha400094c, 32'd17);
pulp_write32(axi_m, 32'ha4000950, 32'd2);
pulp_write32(axi_m, 32'ha4000954, 32'h800019c0);
pulp_write32(axi_m, 32'ha40019c0, 32'h800009d8);
pulp_write32(axi_m, 32'ha40019c4, 32'h80000c94);
pulp_write32(axi_m, 32'ha4000998, 32'h00110000);
pulp_write32(axi_m, 32'ha400099c, 32'h00110001);
pulp_write32(axi_m, 32'ha40009a0, 32'h00110002);
pulp_write32(axi_m, 32'ha40009a4, 32'h00110003);
pulp_write32(axi_m, 32'ha40009a8, 32'h00110004);
pulp_write32(axi_m, 32'ha40009ac, 32'h00110005);
pulp_write32(axi_m, 32'ha40009b0, 32'h00110006);
pulp_write32(axi_m, 32'ha40009b4, 32'h00110007);
pulp_write32(axi_m, 32'ha40009b8, 32'h00110008);
pulp_write32(axi_m, 32'ha40009bc, 32'h00110009);
pulp_write32(axi_m, 32'ha40009c0, 32'h0011000a);
pulp_write32(axi_m, 32'ha40009c4, 32'h0011000b);
pulp_write32(axi_m, 32'ha40009c8, 32'h0011000c);
pulp_write32(axi_m, 32'ha40009cc, 32'h0011000d);
pulp_write32(axi_m, 32'ha40009d0, 32'h0011000e);
pulp_write32(axi_m, 32'ha40009d4, 32'h0011000f);

pulp_write32(axi_m, 32'ha40009d8, 32'd18);
pulp_write32(axi_m, 32'ha40009dc, 32'd1);
pulp_write32(axi_m, 32'ha40009e0, 32'h800019c8);
pulp_write32(axi_m, 32'ha40019c8, 32'h80000d20);
pulp_write32(axi_m, 32'ha4000a24, 32'h00120000);
pulp_write32(axi_m, 32'ha4000a28, 32'h00120001);
pulp_write32(axi_m, 32'ha4000a2c, 32'h00120002);
pulp_write32(axi_m, 32'ha4000a30, 32'h00120003);
pulp_write32(axi_m, 32'ha4000a34, 32'h00120004);
pulp_write32(axi_m, 32'ha4000a38, 32'h00120005);
pulp_write32(axi_m, 32'ha4000a3c, 32'h00120006);
pulp_write32(axi_m, 32'ha4000a40, 32'h00120007);
pulp_write32(axi_m, 32'ha4000a44, 32'h00120008);
pulp_write32(axi_m, 32'ha4000a48, 32'h00120009);
pulp_write32(axi_m, 32'ha4000a4c, 32'h0012000a);
pulp_write32(axi_m, 32'ha4000a50, 32'h0012000b);
pulp_write32(axi_m, 32'ha4000a54, 32'h0012000c);
pulp_write32(axi_m, 32'ha4000a58, 32'h0012000d);
pulp_write32(axi_m, 32'ha4000a5c, 32'h0012000e);
pulp_write32(axi_m, 32'ha4000a60, 32'h0012000f);

pulp_write32(axi_m, 32'ha4000a64, 32'd19);
pulp_write32(axi_m, 32'ha4000a68, 32'd2);
pulp_write32(axi_m, 32'ha4000a6c, 32'h800019d0);
pulp_write32(axi_m, 32'ha40019d0, 32'h80000dac);
pulp_write32(axi_m, 32'ha40019d4, 32'h800015e0);
pulp_write32(axi_m, 32'ha4000ab0, 32'h00130000);
pulp_write32(axi_m, 32'ha4000ab4, 32'h00130001);
pulp_write32(axi_m, 32'ha4000ab8, 32'h00130002);
pulp_write32(axi_m, 32'ha4000abc, 32'h00130003);
pulp_write32(axi_m, 32'ha4000ac0, 32'h00130004);
pulp_write32(axi_m, 32'ha4000ac4, 32'h00130005);
pulp_write32(axi_m, 32'ha4000ac8, 32'h00130006);
pulp_write32(axi_m, 32'ha4000acc, 32'h00130007);
pulp_write32(axi_m, 32'ha4000ad0, 32'h00130008);
pulp_write32(axi_m, 32'ha4000ad4, 32'h00130009);
pulp_write32(axi_m, 32'ha4000ad8, 32'h0013000a);
pulp_write32(axi_m, 32'ha4000adc, 32'h0013000b);
pulp_write32(axi_m, 32'ha4000ae0, 32'h0013000c);
pulp_write32(axi_m, 32'ha4000ae4, 32'h0013000d);
pulp_write32(axi_m, 32'ha4000ae8, 32'h0013000e);
pulp_write32(axi_m, 32'ha4000aec, 32'h0013000f);

pulp_write32(axi_m, 32'ha4000af0, 32'd20);
pulp_write32(axi_m, 32'ha4000af4, 32'd2);
pulp_write32(axi_m, 32'ha4000af8, 32'h800019d8);
pulp_write32(axi_m, 32'ha40019d8, 32'h80000b7c);
pulp_write32(axi_m, 32'ha40019dc, 32'h80000c08);
pulp_write32(axi_m, 32'ha4000b3c, 32'h00140000);
pulp_write32(axi_m, 32'ha4000b40, 32'h00140001);
pulp_write32(axi_m, 32'ha4000b44, 32'h00140002);
pulp_write32(axi_m, 32'ha4000b48, 32'h00140003);
pulp_write32(axi_m, 32'ha4000b4c, 32'h00140004);
pulp_write32(axi_m, 32'ha4000b50, 32'h00140005);
pulp_write32(axi_m, 32'ha4000b54, 32'h00140006);
pulp_write32(axi_m, 32'ha4000b58, 32'h00140007);
pulp_write32(axi_m, 32'ha4000b5c, 32'h00140008);
pulp_write32(axi_m, 32'ha4000b60, 32'h00140009);
pulp_write32(axi_m, 32'ha4000b64, 32'h0014000a);
pulp_write32(axi_m, 32'ha4000b68, 32'h0014000b);
pulp_write32(axi_m, 32'ha4000b6c, 32'h0014000c);
pulp_write32(axi_m, 32'ha4000b70, 32'h0014000d);
pulp_write32(axi_m, 32'ha4000b74, 32'h0014000e);
pulp_write32(axi_m, 32'ha4000b78, 32'h0014000f);

pulp_write32(axi_m, 32'ha4000b7c, 32'd21);
pulp_write32(axi_m, 32'ha4000b80, 32'd0);
pulp_write32(axi_m, 32'ha4000bc8, 32'h00150000);
pulp_write32(axi_m, 32'ha4000bcc, 32'h00150001);
pulp_write32(axi_m, 32'ha4000bd0, 32'h00150002);
pulp_write32(axi_m, 32'ha4000bd4, 32'h00150003);
pulp_write32(axi_m, 32'ha4000bd8, 32'h00150004);
pulp_write32(axi_m, 32'ha4000bdc, 32'h00150005);
pulp_write32(axi_m, 32'ha4000be0, 32'h00150006);
pulp_write32(axi_m, 32'ha4000be4, 32'h00150007);
pulp_write32(axi_m, 32'ha4000be8, 32'h00150008);
pulp_write32(axi_m, 32'ha4000bec, 32'h00150009);
pulp_write32(axi_m, 32'ha4000bf0, 32'h0015000a);
pulp_write32(axi_m, 32'ha4000bf4, 32'h0015000b);
pulp_write32(axi_m, 32'ha4000bf8, 32'h0015000c);
pulp_write32(axi_m, 32'ha4000bfc, 32'h0015000d);
pulp_write32(axi_m, 32'ha4000c00, 32'h0015000e);
pulp_write32(axi_m, 32'ha4000c04, 32'h0015000f);

pulp_write32(axi_m, 32'ha4000c08, 32'd22);
pulp_write32(axi_m, 32'ha4000c0c, 32'd1);
pulp_write32(axi_m, 32'ha4000c10, 32'h800019e0);
pulp_write32(axi_m, 32'ha40019e0, 32'h80000c94);
pulp_write32(axi_m, 32'ha4000c54, 32'h00160000);
pulp_write32(axi_m, 32'ha4000c58, 32'h00160001);
pulp_write32(axi_m, 32'ha4000c5c, 32'h00160002);
pulp_write32(axi_m, 32'ha4000c60, 32'h00160003);
pulp_write32(axi_m, 32'ha4000c64, 32'h00160004);
pulp_write32(axi_m, 32'ha4000c68, 32'h00160005);
pulp_write32(axi_m, 32'ha4000c6c, 32'h00160006);
pulp_write32(axi_m, 32'ha4000c70, 32'h00160007);
pulp_write32(axi_m, 32'ha4000c74, 32'h00160008);
pulp_write32(axi_m, 32'ha4000c78, 32'h00160009);
pulp_write32(axi_m, 32'ha4000c7c, 32'h0016000a);
pulp_write32(axi_m, 32'ha4000c80, 32'h0016000b);
pulp_write32(axi_m, 32'ha4000c84, 32'h0016000c);
pulp_write32(axi_m, 32'ha4000c88, 32'h0016000d);
pulp_write32(axi_m, 32'ha4000c8c, 32'h0016000e);
pulp_write32(axi_m, 32'ha4000c90, 32'h0016000f);

pulp_write32(axi_m, 32'ha4000c94, 32'd23);
pulp_write32(axi_m, 32'ha4000c98, 32'd1);
pulp_write32(axi_m, 32'ha4000c9c, 32'h800019e8);
pulp_write32(axi_m, 32'ha40019e8, 32'h80000d20);
pulp_write32(axi_m, 32'ha4000ce0, 32'h00170000);
pulp_write32(axi_m, 32'ha4000ce4, 32'h00170001);
pulp_write32(axi_m, 32'ha4000ce8, 32'h00170002);
pulp_write32(axi_m, 32'ha4000cec, 32'h00170003);
pulp_write32(axi_m, 32'ha4000cf0, 32'h00170004);
pulp_write32(axi_m, 32'ha4000cf4, 32'h00170005);
pulp_write32(axi_m, 32'ha4000cf8, 32'h00170006);
pulp_write32(axi_m, 32'ha4000cfc, 32'h00170007);
pulp_write32(axi_m, 32'ha4000d00, 32'h00170008);
pulp_write32(axi_m, 32'ha4000d04, 32'h00170009);
pulp_write32(axi_m, 32'ha4000d08, 32'h0017000a);
pulp_write32(axi_m, 32'ha4000d0c, 32'h0017000b);
pulp_write32(axi_m, 32'ha4000d10, 32'h0017000c);
pulp_write32(axi_m, 32'ha4000d14, 32'h0017000d);
pulp_write32(axi_m, 32'ha4000d18, 32'h0017000e);
pulp_write32(axi_m, 32'ha4000d1c, 32'h0017000f);

pulp_write32(axi_m, 32'ha4000d20, 32'd24);
pulp_write32(axi_m, 32'ha4000d24, 32'd0);
pulp_write32(axi_m, 32'ha4000d6c, 32'h00180000);
pulp_write32(axi_m, 32'ha4000d70, 32'h00180001);
pulp_write32(axi_m, 32'ha4000d74, 32'h00180002);
pulp_write32(axi_m, 32'ha4000d78, 32'h00180003);
pulp_write32(axi_m, 32'ha4000d7c, 32'h00180004);
pulp_write32(axi_m, 32'ha4000d80, 32'h00180005);
pulp_write32(axi_m, 32'ha4000d84, 32'h00180006);
pulp_write32(axi_m, 32'ha4000d88, 32'h00180007);
pulp_write32(axi_m, 32'ha4000d8c, 32'h00180008);
pulp_write32(axi_m, 32'ha4000d90, 32'h00180009);
pulp_write32(axi_m, 32'ha4000d94, 32'h0018000a);
pulp_write32(axi_m, 32'ha4000d98, 32'h0018000b);
pulp_write32(axi_m, 32'ha4000d9c, 32'h0018000c);
pulp_write32(axi_m, 32'ha4000da0, 32'h0018000d);
pulp_write32(axi_m, 32'ha4000da4, 32'h0018000e);
pulp_write32(axi_m, 32'ha4000da8, 32'h0018000f);

pulp_write32(axi_m, 32'ha4000dac, 32'd25);
pulp_write32(axi_m, 32'ha4000db0, 32'd2);
pulp_write32(axi_m, 32'ha4000db4, 32'h800019f0);
pulp_write32(axi_m, 32'ha40019f0, 32'h80000e38);
pulp_write32(axi_m, 32'ha40019f4, 32'h800014c8);
pulp_write32(axi_m, 32'ha4000df8, 32'h00190000);
pulp_write32(axi_m, 32'ha4000dfc, 32'h00190001);
pulp_write32(axi_m, 32'ha4000e00, 32'h00190002);
pulp_write32(axi_m, 32'ha4000e04, 32'h00190003);
pulp_write32(axi_m, 32'ha4000e08, 32'h00190004);
pulp_write32(axi_m, 32'ha4000e0c, 32'h00190005);
pulp_write32(axi_m, 32'ha4000e10, 32'h00190006);
pulp_write32(axi_m, 32'ha4000e14, 32'h00190007);
pulp_write32(axi_m, 32'ha4000e18, 32'h00190008);
pulp_write32(axi_m, 32'ha4000e1c, 32'h00190009);
pulp_write32(axi_m, 32'ha4000e20, 32'h0019000a);
pulp_write32(axi_m, 32'ha4000e24, 32'h0019000b);
pulp_write32(axi_m, 32'ha4000e28, 32'h0019000c);
pulp_write32(axi_m, 32'ha4000e2c, 32'h0019000d);
pulp_write32(axi_m, 32'ha4000e30, 32'h0019000e);
pulp_write32(axi_m, 32'ha4000e34, 32'h0019000f);

pulp_write32(axi_m, 32'ha4000e38, 32'd26);
pulp_write32(axi_m, 32'ha4000e3c, 32'd1);
pulp_write32(axi_m, 32'ha4000e40, 32'h800019f8);
pulp_write32(axi_m, 32'ha40019f8, 32'h80001298);
pulp_write32(axi_m, 32'ha4000e84, 32'h001a0000);
pulp_write32(axi_m, 32'ha4000e88, 32'h001a0001);
pulp_write32(axi_m, 32'ha4000e8c, 32'h001a0002);
pulp_write32(axi_m, 32'ha4000e90, 32'h001a0003);
pulp_write32(axi_m, 32'ha4000e94, 32'h001a0004);
pulp_write32(axi_m, 32'ha4000e98, 32'h001a0005);
pulp_write32(axi_m, 32'ha4000e9c, 32'h001a0006);
pulp_write32(axi_m, 32'ha4000ea0, 32'h001a0007);
pulp_write32(axi_m, 32'ha4000ea4, 32'h001a0008);
pulp_write32(axi_m, 32'ha4000ea8, 32'h001a0009);
pulp_write32(axi_m, 32'ha4000eac, 32'h001a000a);
pulp_write32(axi_m, 32'ha4000eb0, 32'h001a000b);
pulp_write32(axi_m, 32'ha4000eb4, 32'h001a000c);
pulp_write32(axi_m, 32'ha4000eb8, 32'h001a000d);
pulp_write32(axi_m, 32'ha4000ebc, 32'h001a000e);
pulp_write32(axi_m, 32'ha4000ec0, 32'h001a000f);

pulp_write32(axi_m, 32'ha4000ec4, 32'd27);
pulp_write32(axi_m, 32'ha4000ec8, 32'd2);
pulp_write32(axi_m, 32'ha4000ecc, 32'h80001a00);
pulp_write32(axi_m, 32'ha4001a00, 32'h80000f50);
pulp_write32(axi_m, 32'ha4001a04, 32'h80001554);
pulp_write32(axi_m, 32'ha4000f10, 32'h001b0000);
pulp_write32(axi_m, 32'ha4000f14, 32'h001b0001);
pulp_write32(axi_m, 32'ha4000f18, 32'h001b0002);
pulp_write32(axi_m, 32'ha4000f1c, 32'h001b0003);
pulp_write32(axi_m, 32'ha4000f20, 32'h001b0004);
pulp_write32(axi_m, 32'ha4000f24, 32'h001b0005);
pulp_write32(axi_m, 32'ha4000f28, 32'h001b0006);
pulp_write32(axi_m, 32'ha4000f2c, 32'h001b0007);
pulp_write32(axi_m, 32'ha4000f30, 32'h001b0008);
pulp_write32(axi_m, 32'ha4000f34, 32'h001b0009);
pulp_write32(axi_m, 32'ha4000f38, 32'h001b000a);
pulp_write32(axi_m, 32'ha4000f3c, 32'h001b000b);
pulp_write32(axi_m, 32'ha4000f40, 32'h001b000c);
pulp_write32(axi_m, 32'ha4000f44, 32'h001b000d);
pulp_write32(axi_m, 32'ha4000f48, 32'h001b000e);
pulp_write32(axi_m, 32'ha4000f4c, 32'h001b000f);

pulp_write32(axi_m, 32'ha4000f50, 32'd28);
pulp_write32(axi_m, 32'ha4000f54, 32'd1);
pulp_write32(axi_m, 32'ha4000f58, 32'h80001a08);
pulp_write32(axi_m, 32'ha4001a08, 32'h80001298);
pulp_write32(axi_m, 32'ha4000f9c, 32'h001c0000);
pulp_write32(axi_m, 32'ha4000fa0, 32'h001c0001);
pulp_write32(axi_m, 32'ha4000fa4, 32'h001c0002);
pulp_write32(axi_m, 32'ha4000fa8, 32'h001c0003);
pulp_write32(axi_m, 32'ha4000fac, 32'h001c0004);
pulp_write32(axi_m, 32'ha4000fb0, 32'h001c0005);
pulp_write32(axi_m, 32'ha4000fb4, 32'h001c0006);
pulp_write32(axi_m, 32'ha4000fb8, 32'h001c0007);
pulp_write32(axi_m, 32'ha4000fbc, 32'h001c0008);
pulp_write32(axi_m, 32'ha4000fc0, 32'h001c0009);
pulp_write32(axi_m, 32'ha4000fc4, 32'h001c000a);
pulp_write32(axi_m, 32'ha4000fc8, 32'h001c000b);
pulp_write32(axi_m, 32'ha4000fcc, 32'h001c000c);
pulp_write32(axi_m, 32'ha4000fd0, 32'h001c000d);
pulp_write32(axi_m, 32'ha4000fd4, 32'h001c000e);
pulp_write32(axi_m, 32'ha4000fd8, 32'h001c000f);

pulp_write32(axi_m, 32'ha4000fdc, 32'd29);
pulp_write32(axi_m, 32'ha4000fe0, 32'd2);
pulp_write32(axi_m, 32'ha4000fe4, 32'h80001a10);
pulp_write32(axi_m, 32'ha4001a10, 32'h80001068);
pulp_write32(axi_m, 32'ha4001a14, 32'h80001810);
pulp_write32(axi_m, 32'ha4001028, 32'h001d0000);
pulp_write32(axi_m, 32'ha400102c, 32'h001d0001);
pulp_write32(axi_m, 32'ha4001030, 32'h001d0002);
pulp_write32(axi_m, 32'ha4001034, 32'h001d0003);
pulp_write32(axi_m, 32'ha4001038, 32'h001d0004);
pulp_write32(axi_m, 32'ha400103c, 32'h001d0005);
pulp_write32(axi_m, 32'ha4001040, 32'h001d0006);
pulp_write32(axi_m, 32'ha4001044, 32'h001d0007);
pulp_write32(axi_m, 32'ha4001048, 32'h001d0008);
pulp_write32(axi_m, 32'ha400104c, 32'h001d0009);
pulp_write32(axi_m, 32'ha4001050, 32'h001d000a);
pulp_write32(axi_m, 32'ha4001054, 32'h001d000b);
pulp_write32(axi_m, 32'ha4001058, 32'h001d000c);
pulp_write32(axi_m, 32'ha400105c, 32'h001d000d);
pulp_write32(axi_m, 32'ha4001060, 32'h001d000e);
pulp_write32(axi_m, 32'ha4001064, 32'h001d000f);

pulp_write32(axi_m, 32'ha4001068, 32'd30);
pulp_write32(axi_m, 32'ha400106c, 32'd1);
pulp_write32(axi_m, 32'ha4001070, 32'h80001a18);
pulp_write32(axi_m, 32'ha4001a18, 32'h80001324);
pulp_write32(axi_m, 32'ha40010b4, 32'h001e0000);
pulp_write32(axi_m, 32'ha40010b8, 32'h001e0001);
pulp_write32(axi_m, 32'ha40010bc, 32'h001e0002);
pulp_write32(axi_m, 32'ha40010c0, 32'h001e0003);
pulp_write32(axi_m, 32'ha40010c4, 32'h001e0004);
pulp_write32(axi_m, 32'ha40010c8, 32'h001e0005);
pulp_write32(axi_m, 32'ha40010cc, 32'h001e0006);
pulp_write32(axi_m, 32'ha40010d0, 32'h001e0007);
pulp_write32(axi_m, 32'ha40010d4, 32'h001e0008);
pulp_write32(axi_m, 32'ha40010d8, 32'h001e0009);
pulp_write32(axi_m, 32'ha40010dc, 32'h001e000a);
pulp_write32(axi_m, 32'ha40010e0, 32'h001e000b);
pulp_write32(axi_m, 32'ha40010e4, 32'h001e000c);
pulp_write32(axi_m, 32'ha40010e8, 32'h001e000d);
pulp_write32(axi_m, 32'ha40010ec, 32'h001e000e);
pulp_write32(axi_m, 32'ha40010f0, 32'h001e000f);

pulp_write32(axi_m, 32'ha40010f4, 32'd31);
pulp_write32(axi_m, 32'ha40010f8, 32'd2);
pulp_write32(axi_m, 32'ha40010fc, 32'h80001a20);
pulp_write32(axi_m, 32'ha4001a20, 32'h80001180);
pulp_write32(axi_m, 32'ha4001a24, 32'h80001324);
pulp_write32(axi_m, 32'ha4001140, 32'h001f0000);
pulp_write32(axi_m, 32'ha4001144, 32'h001f0001);
pulp_write32(axi_m, 32'ha4001148, 32'h001f0002);
pulp_write32(axi_m, 32'ha400114c, 32'h001f0003);
pulp_write32(axi_m, 32'ha4001150, 32'h001f0004);
pulp_write32(axi_m, 32'ha4001154, 32'h001f0005);
pulp_write32(axi_m, 32'ha4001158, 32'h001f0006);
pulp_write32(axi_m, 32'ha400115c, 32'h001f0007);
pulp_write32(axi_m, 32'ha4001160, 32'h001f0008);
pulp_write32(axi_m, 32'ha4001164, 32'h001f0009);
pulp_write32(axi_m, 32'ha4001168, 32'h001f000a);
pulp_write32(axi_m, 32'ha400116c, 32'h001f000b);
pulp_write32(axi_m, 32'ha4001170, 32'h001f000c);
pulp_write32(axi_m, 32'ha4001174, 32'h001f000d);
pulp_write32(axi_m, 32'ha4001178, 32'h001f000e);
pulp_write32(axi_m, 32'ha400117c, 32'h001f000f);

pulp_write32(axi_m, 32'ha4001180, 32'd32);
pulp_write32(axi_m, 32'ha4001184, 32'd2);
pulp_write32(axi_m, 32'ha4001188, 32'h80001a28);
pulp_write32(axi_m, 32'ha4001a28, 32'h8000120c);
pulp_write32(axi_m, 32'ha4001a2c, 32'h800016f8);
pulp_write32(axi_m, 32'ha40011cc, 32'h00200000);
pulp_write32(axi_m, 32'ha40011d0, 32'h00200001);
pulp_write32(axi_m, 32'ha40011d4, 32'h00200002);
pulp_write32(axi_m, 32'ha40011d8, 32'h00200003);
pulp_write32(axi_m, 32'ha40011dc, 32'h00200004);
pulp_write32(axi_m, 32'ha40011e0, 32'h00200005);
pulp_write32(axi_m, 32'ha40011e4, 32'h00200006);
pulp_write32(axi_m, 32'ha40011e8, 32'h00200007);
pulp_write32(axi_m, 32'ha40011ec, 32'h00200008);
pulp_write32(axi_m, 32'ha40011f0, 32'h00200009);
pulp_write32(axi_m, 32'ha40011f4, 32'h0020000a);
pulp_write32(axi_m, 32'ha40011f8, 32'h0020000b);
pulp_write32(axi_m, 32'ha40011fc, 32'h0020000c);
pulp_write32(axi_m, 32'ha4001200, 32'h0020000d);
pulp_write32(axi_m, 32'ha4001204, 32'h0020000e);
pulp_write32(axi_m, 32'ha4001208, 32'h0020000f);

pulp_write32(axi_m, 32'ha400120c, 32'd33);
pulp_write32(axi_m, 32'ha4001210, 32'd1);
pulp_write32(axi_m, 32'ha4001214, 32'h80001a30);
pulp_write32(axi_m, 32'ha4001a30, 32'h80001784);
pulp_write32(axi_m, 32'ha4001258, 32'h00210000);
pulp_write32(axi_m, 32'ha400125c, 32'h00210001);
pulp_write32(axi_m, 32'ha4001260, 32'h00210002);
pulp_write32(axi_m, 32'ha4001264, 32'h00210003);
pulp_write32(axi_m, 32'ha4001268, 32'h00210004);
pulp_write32(axi_m, 32'ha400126c, 32'h00210005);
pulp_write32(axi_m, 32'ha4001270, 32'h00210006);
pulp_write32(axi_m, 32'ha4001274, 32'h00210007);
pulp_write32(axi_m, 32'ha4001278, 32'h00210008);
pulp_write32(axi_m, 32'ha400127c, 32'h00210009);
pulp_write32(axi_m, 32'ha4001280, 32'h0021000a);
pulp_write32(axi_m, 32'ha4001284, 32'h0021000b);
pulp_write32(axi_m, 32'ha4001288, 32'h0021000c);
pulp_write32(axi_m, 32'ha400128c, 32'h0021000d);
pulp_write32(axi_m, 32'ha4001290, 32'h0021000e);
pulp_write32(axi_m, 32'ha4001294, 32'h0021000f);

pulp_write32(axi_m, 32'ha4001298, 32'd34);
pulp_write32(axi_m, 32'ha400129c, 32'd1);
pulp_write32(axi_m, 32'ha40012a0, 32'h80001a38);
pulp_write32(axi_m, 32'ha4001a38, 32'h800013b0);
pulp_write32(axi_m, 32'ha40012e4, 32'h00220000);
pulp_write32(axi_m, 32'ha40012e8, 32'h00220001);
pulp_write32(axi_m, 32'ha40012ec, 32'h00220002);
pulp_write32(axi_m, 32'ha40012f0, 32'h00220003);
pulp_write32(axi_m, 32'ha40012f4, 32'h00220004);
pulp_write32(axi_m, 32'ha40012f8, 32'h00220005);
pulp_write32(axi_m, 32'ha40012fc, 32'h00220006);
pulp_write32(axi_m, 32'ha4001300, 32'h00220007);
pulp_write32(axi_m, 32'ha4001304, 32'h00220008);
pulp_write32(axi_m, 32'ha4001308, 32'h00220009);
pulp_write32(axi_m, 32'ha400130c, 32'h0022000a);
pulp_write32(axi_m, 32'ha4001310, 32'h0022000b);
pulp_write32(axi_m, 32'ha4001314, 32'h0022000c);
pulp_write32(axi_m, 32'ha4001318, 32'h0022000d);
pulp_write32(axi_m, 32'ha400131c, 32'h0022000e);
pulp_write32(axi_m, 32'ha4001320, 32'h0022000f);

pulp_write32(axi_m, 32'ha4001324, 32'd35);
pulp_write32(axi_m, 32'ha4001328, 32'd1);
pulp_write32(axi_m, 32'ha400132c, 32'h80001a40);
pulp_write32(axi_m, 32'ha4001a40, 32'h8000143c);
pulp_write32(axi_m, 32'ha4001370, 32'h00230000);
pulp_write32(axi_m, 32'ha4001374, 32'h00230001);
pulp_write32(axi_m, 32'ha4001378, 32'h00230002);
pulp_write32(axi_m, 32'ha400137c, 32'h00230003);
pulp_write32(axi_m, 32'ha4001380, 32'h00230004);
pulp_write32(axi_m, 32'ha4001384, 32'h00230005);
pulp_write32(axi_m, 32'ha4001388, 32'h00230006);
pulp_write32(axi_m, 32'ha400138c, 32'h00230007);
pulp_write32(axi_m, 32'ha4001390, 32'h00230008);
pulp_write32(axi_m, 32'ha4001394, 32'h00230009);
pulp_write32(axi_m, 32'ha4001398, 32'h0023000a);
pulp_write32(axi_m, 32'ha400139c, 32'h0023000b);
pulp_write32(axi_m, 32'ha40013a0, 32'h0023000c);
pulp_write32(axi_m, 32'ha40013a4, 32'h0023000d);
pulp_write32(axi_m, 32'ha40013a8, 32'h0023000e);
pulp_write32(axi_m, 32'ha40013ac, 32'h0023000f);

pulp_write32(axi_m, 32'ha40013b0, 32'd36);
pulp_write32(axi_m, 32'ha40013b4, 32'd2);
pulp_write32(axi_m, 32'ha40013b8, 32'h80001a48);
pulp_write32(axi_m, 32'ha4001a48, 32'h800014c8);
pulp_write32(axi_m, 32'ha4001a4c, 32'h80001554);
pulp_write32(axi_m, 32'ha40013fc, 32'h00240000);
pulp_write32(axi_m, 32'ha4001400, 32'h00240001);
pulp_write32(axi_m, 32'ha4001404, 32'h00240002);
pulp_write32(axi_m, 32'ha4001408, 32'h00240003);
pulp_write32(axi_m, 32'ha400140c, 32'h00240004);
pulp_write32(axi_m, 32'ha4001410, 32'h00240005);
pulp_write32(axi_m, 32'ha4001414, 32'h00240006);
pulp_write32(axi_m, 32'ha4001418, 32'h00240007);
pulp_write32(axi_m, 32'ha400141c, 32'h00240008);
pulp_write32(axi_m, 32'ha4001420, 32'h00240009);
pulp_write32(axi_m, 32'ha4001424, 32'h0024000a);
pulp_write32(axi_m, 32'ha4001428, 32'h0024000b);
pulp_write32(axi_m, 32'ha400142c, 32'h0024000c);
pulp_write32(axi_m, 32'ha4001430, 32'h0024000d);
pulp_write32(axi_m, 32'ha4001434, 32'h0024000e);
pulp_write32(axi_m, 32'ha4001438, 32'h0024000f);

pulp_write32(axi_m, 32'ha400143c, 32'd37);
pulp_write32(axi_m, 32'ha4001440, 32'd2);
pulp_write32(axi_m, 32'ha4001444, 32'h80001a50);
pulp_write32(axi_m, 32'ha4001a50, 32'h800016f8);
pulp_write32(axi_m, 32'ha4001a54, 32'h80001810);
pulp_write32(axi_m, 32'ha4001488, 32'h00250000);
pulp_write32(axi_m, 32'ha400148c, 32'h00250001);
pulp_write32(axi_m, 32'ha4001490, 32'h00250002);
pulp_write32(axi_m, 32'ha4001494, 32'h00250003);
pulp_write32(axi_m, 32'ha4001498, 32'h00250004);
pulp_write32(axi_m, 32'ha400149c, 32'h00250005);
pulp_write32(axi_m, 32'ha40014a0, 32'h00250006);
pulp_write32(axi_m, 32'ha40014a4, 32'h00250007);
pulp_write32(axi_m, 32'ha40014a8, 32'h00250008);
pulp_write32(axi_m, 32'ha40014ac, 32'h00250009);
pulp_write32(axi_m, 32'ha40014b0, 32'h0025000a);
pulp_write32(axi_m, 32'ha40014b4, 32'h0025000b);
pulp_write32(axi_m, 32'ha40014b8, 32'h0025000c);
pulp_write32(axi_m, 32'ha40014bc, 32'h0025000d);
pulp_write32(axi_m, 32'ha40014c0, 32'h0025000e);
pulp_write32(axi_m, 32'ha40014c4, 32'h0025000f);

pulp_write32(axi_m, 32'ha40014c8, 32'd38);
pulp_write32(axi_m, 32'ha40014cc, 32'd1);
pulp_write32(axi_m, 32'ha40014d0, 32'h80001a58);
pulp_write32(axi_m, 32'ha4001a58, 32'h800015e0);
pulp_write32(axi_m, 32'ha4001514, 32'h00260000);
pulp_write32(axi_m, 32'ha4001518, 32'h00260001);
pulp_write32(axi_m, 32'ha400151c, 32'h00260002);
pulp_write32(axi_m, 32'ha4001520, 32'h00260003);
pulp_write32(axi_m, 32'ha4001524, 32'h00260004);
pulp_write32(axi_m, 32'ha4001528, 32'h00260005);
pulp_write32(axi_m, 32'ha400152c, 32'h00260006);
pulp_write32(axi_m, 32'ha4001530, 32'h00260007);
pulp_write32(axi_m, 32'ha4001534, 32'h00260008);
pulp_write32(axi_m, 32'ha4001538, 32'h00260009);
pulp_write32(axi_m, 32'ha400153c, 32'h0026000a);
pulp_write32(axi_m, 32'ha4001540, 32'h0026000b);
pulp_write32(axi_m, 32'ha4001544, 32'h0026000c);
pulp_write32(axi_m, 32'ha4001548, 32'h0026000d);
pulp_write32(axi_m, 32'ha400154c, 32'h0026000e);
pulp_write32(axi_m, 32'ha4001550, 32'h0026000f);

pulp_write32(axi_m, 32'ha4001554, 32'd39);
pulp_write32(axi_m, 32'ha4001558, 32'd1);
pulp_write32(axi_m, 32'ha400155c, 32'h80001a60);
pulp_write32(axi_m, 32'ha4001a60, 32'h8000166c);
pulp_write32(axi_m, 32'ha40015a0, 32'h00270000);
pulp_write32(axi_m, 32'ha40015a4, 32'h00270001);
pulp_write32(axi_m, 32'ha40015a8, 32'h00270002);
pulp_write32(axi_m, 32'ha40015ac, 32'h00270003);
pulp_write32(axi_m, 32'ha40015b0, 32'h00270004);
pulp_write32(axi_m, 32'ha40015b4, 32'h00270005);
pulp_write32(axi_m, 32'ha40015b8, 32'h00270006);
pulp_write32(axi_m, 32'ha40015bc, 32'h00270007);
pulp_write32(axi_m, 32'ha40015c0, 32'h00270008);
pulp_write32(axi_m, 32'ha40015c4, 32'h00270009);
pulp_write32(axi_m, 32'ha40015c8, 32'h0027000a);
pulp_write32(axi_m, 32'ha40015cc, 32'h0027000b);
pulp_write32(axi_m, 32'ha40015d0, 32'h0027000c);
pulp_write32(axi_m, 32'ha40015d4, 32'h0027000d);
pulp_write32(axi_m, 32'ha40015d8, 32'h0027000e);
pulp_write32(axi_m, 32'ha40015dc, 32'h0027000f);

pulp_write32(axi_m, 32'ha40015e0, 32'd40);
pulp_write32(axi_m, 32'ha40015e4, 32'd1);
pulp_write32(axi_m, 32'ha40015e8, 32'h80001a68);
pulp_write32(axi_m, 32'ha4001a68, 32'h8000166c);
pulp_write32(axi_m, 32'ha400162c, 32'h00280000);
pulp_write32(axi_m, 32'ha4001630, 32'h00280001);
pulp_write32(axi_m, 32'ha4001634, 32'h00280002);
pulp_write32(axi_m, 32'ha4001638, 32'h00280003);
pulp_write32(axi_m, 32'ha400163c, 32'h00280004);
pulp_write32(axi_m, 32'ha4001640, 32'h00280005);
pulp_write32(axi_m, 32'ha4001644, 32'h00280006);
pulp_write32(axi_m, 32'ha4001648, 32'h00280007);
pulp_write32(axi_m, 32'ha400164c, 32'h00280008);
pulp_write32(axi_m, 32'ha4001650, 32'h00280009);
pulp_write32(axi_m, 32'ha4001654, 32'h0028000a);
pulp_write32(axi_m, 32'ha4001658, 32'h0028000b);
pulp_write32(axi_m, 32'ha400165c, 32'h0028000c);
pulp_write32(axi_m, 32'ha4001660, 32'h0028000d);
pulp_write32(axi_m, 32'ha4001664, 32'h0028000e);
pulp_write32(axi_m, 32'ha4001668, 32'h0028000f);

pulp_write32(axi_m, 32'ha400166c, 32'd41);
pulp_write32(axi_m, 32'ha4001670, 32'd0);
pulp_write32(axi_m, 32'ha40016b8, 32'h00290000);
pulp_write32(axi_m, 32'ha40016bc, 32'h00290001);
pulp_write32(axi_m, 32'ha40016c0, 32'h00290002);
pulp_write32(axi_m, 32'ha40016c4, 32'h00290003);
pulp_write32(axi_m, 32'ha40016c8, 32'h00290004);
pulp_write32(axi_m, 32'ha40016cc, 32'h00290005);
pulp_write32(axi_m, 32'ha40016d0, 32'h00290006);
pulp_write32(axi_m, 32'ha40016d4, 32'h00290007);
pulp_write32(axi_m, 32'ha40016d8, 32'h00290008);
pulp_write32(axi_m, 32'ha40016dc, 32'h00290009);
pulp_write32(axi_m, 32'ha40016e0, 32'h0029000a);
pulp_write32(axi_m, 32'ha40016e4, 32'h0029000b);
pulp_write32(axi_m, 32'ha40016e8, 32'h0029000c);
pulp_write32(axi_m, 32'ha40016ec, 32'h0029000d);
pulp_write32(axi_m, 32'ha40016f0, 32'h0029000e);
pulp_write32(axi_m, 32'ha40016f4, 32'h0029000f);

pulp_write32(axi_m, 32'ha40016f8, 32'd42);
pulp_write32(axi_m, 32'ha40016fc, 32'd1);
pulp_write32(axi_m, 32'ha4001700, 32'h80001a70);
pulp_write32(axi_m, 32'ha4001a70, 32'h80001784);
pulp_write32(axi_m, 32'ha4001744, 32'h002a0000);
pulp_write32(axi_m, 32'ha4001748, 32'h002a0001);
pulp_write32(axi_m, 32'ha400174c, 32'h002a0002);
pulp_write32(axi_m, 32'ha4001750, 32'h002a0003);
pulp_write32(axi_m, 32'ha4001754, 32'h002a0004);
pulp_write32(axi_m, 32'ha4001758, 32'h002a0005);
pulp_write32(axi_m, 32'ha400175c, 32'h002a0006);
pulp_write32(axi_m, 32'ha4001760, 32'h002a0007);
pulp_write32(axi_m, 32'ha4001764, 32'h002a0008);
pulp_write32(axi_m, 32'ha4001768, 32'h002a0009);
pulp_write32(axi_m, 32'ha400176c, 32'h002a000a);
pulp_write32(axi_m, 32'ha4001770, 32'h002a000b);
pulp_write32(axi_m, 32'ha4001774, 32'h002a000c);
pulp_write32(axi_m, 32'ha4001778, 32'h002a000d);
pulp_write32(axi_m, 32'ha400177c, 32'h002a000e);
pulp_write32(axi_m, 32'ha4001780, 32'h002a000f);

pulp_write32(axi_m, 32'ha4001784, 32'd43);
pulp_write32(axi_m, 32'ha4001788, 32'd1);
pulp_write32(axi_m, 32'ha400178c, 32'h80001a78);
pulp_write32(axi_m, 32'ha4001a78, 32'h8000189c);
pulp_write32(axi_m, 32'ha40017d0, 32'h002b0000);
pulp_write32(axi_m, 32'ha40017d4, 32'h002b0001);
pulp_write32(axi_m, 32'ha40017d8, 32'h002b0002);
pulp_write32(axi_m, 32'ha40017dc, 32'h002b0003);
pulp_write32(axi_m, 32'ha40017e0, 32'h002b0004);
pulp_write32(axi_m, 32'ha40017e4, 32'h002b0005);
pulp_write32(axi_m, 32'ha40017e8, 32'h002b0006);
pulp_write32(axi_m, 32'ha40017ec, 32'h002b0007);
pulp_write32(axi_m, 32'ha40017f0, 32'h002b0008);
pulp_write32(axi_m, 32'ha40017f4, 32'h002b0009);
pulp_write32(axi_m, 32'ha40017f8, 32'h002b000a);
pulp_write32(axi_m, 32'ha40017fc, 32'h002b000b);
pulp_write32(axi_m, 32'ha4001800, 32'h002b000c);
pulp_write32(axi_m, 32'ha4001804, 32'h002b000d);
pulp_write32(axi_m, 32'ha4001808, 32'h002b000e);
pulp_write32(axi_m, 32'ha400180c, 32'h002b000f);

pulp_write32(axi_m, 32'ha4001810, 32'd44);
pulp_write32(axi_m, 32'ha4001814, 32'd1);
pulp_write32(axi_m, 32'ha4001818, 32'h80001a80);
pulp_write32(axi_m, 32'ha4001a80, 32'h8000189c);
pulp_write32(axi_m, 32'ha400185c, 32'h002c0000);
pulp_write32(axi_m, 32'ha4001860, 32'h002c0001);
pulp_write32(axi_m, 32'ha4001864, 32'h002c0002);
pulp_write32(axi_m, 32'ha4001868, 32'h002c0003);
pulp_write32(axi_m, 32'ha400186c, 32'h002c0004);
pulp_write32(axi_m, 32'ha4001870, 32'h002c0005);
pulp_write32(axi_m, 32'ha4001874, 32'h002c0006);
pulp_write32(axi_m, 32'ha4001878, 32'h002c0007);
pulp_write32(axi_m, 32'ha400187c, 32'h002c0008);
pulp_write32(axi_m, 32'ha4001880, 32'h002c0009);
pulp_write32(axi_m, 32'ha4001884, 32'h002c000a);
pulp_write32(axi_m, 32'ha4001888, 32'h002c000b);
pulp_write32(axi_m, 32'ha400188c, 32'h002c000c);
pulp_write32(axi_m, 32'ha4001890, 32'h002c000d);
pulp_write32(axi_m, 32'ha4001894, 32'h002c000e);
pulp_write32(axi_m, 32'ha4001898, 32'h002c000f);

pulp_write32(axi_m, 32'ha400189c, 32'd45);
pulp_write32(axi_m, 32'ha40018a0, 32'd0);
pulp_write32(axi_m, 32'ha40018e8, 32'h002d0000);
pulp_write32(axi_m, 32'ha40018ec, 32'h002d0001);
pulp_write32(axi_m, 32'ha40018f0, 32'h002d0002);
pulp_write32(axi_m, 32'ha40018f4, 32'h002d0003);
pulp_write32(axi_m, 32'ha40018f8, 32'h002d0004);
pulp_write32(axi_m, 32'ha40018fc, 32'h002d0005);
pulp_write32(axi_m, 32'ha4001900, 32'h002d0006);
pulp_write32(axi_m, 32'ha4001904, 32'h002d0007);
pulp_write32(axi_m, 32'ha4001908, 32'h002d0008);
pulp_write32(axi_m, 32'ha400190c, 32'h002d0009);
pulp_write32(axi_m, 32'ha4001910, 32'h002d000a);
pulp_write32(axi_m, 32'ha4001914, 32'h002d000b);
pulp_write32(axi_m, 32'ha4001918, 32'h002d000c);
pulp_write32(axi_m, 32'ha400191c, 32'h002d000d);
pulp_write32(axi_m, 32'ha4001920, 32'h002d000e);
pulp_write32(axi_m, 32'ha4001924, 32'h002d000f);

