pulp_write32(axi_m, 32'h66000000, 32'd0);
pulp_write32(axi_m, 32'h66000004, 32'd3);
pulp_write32(axi_m, 32'h66000008, 32'h80001928);
pulp_write32(axi_m, 32'h66001928, 32'h80000578);
pulp_write32(axi_m, 32'h6600192c, 32'h80000604);
pulp_write32(axi_m, 32'h66001930, 32'h80000690);
pulp_write32(axi_m, 32'h6600004c, 32'h00000000);
pulp_write32(axi_m, 32'h66000050, 32'h00000001);
pulp_write32(axi_m, 32'h66000054, 32'h00000002);
pulp_write32(axi_m, 32'h66000058, 32'h00000003);
pulp_write32(axi_m, 32'h6600005c, 32'h00000004);
pulp_write32(axi_m, 32'h66000060, 32'h00000005);
pulp_write32(axi_m, 32'h66000064, 32'h00000006);
pulp_write32(axi_m, 32'h66000068, 32'h00000007);
pulp_write32(axi_m, 32'h6600006c, 32'h00000008);
pulp_write32(axi_m, 32'h66000070, 32'h00000009);
pulp_write32(axi_m, 32'h66000074, 32'h0000000a);
pulp_write32(axi_m, 32'h66000078, 32'h0000000b);
pulp_write32(axi_m, 32'h6600007c, 32'h0000000c);
pulp_write32(axi_m, 32'h66000080, 32'h0000000d);
pulp_write32(axi_m, 32'h66000084, 32'h0000000e);
pulp_write32(axi_m, 32'h66000088, 32'h0000000f);

pulp_write32(axi_m, 32'h6600008c, 32'd1);
pulp_write32(axi_m, 32'h66000090, 32'd3);
pulp_write32(axi_m, 32'h66000094, 32'h80001938);
pulp_write32(axi_m, 32'h66001938, 32'h80000118);
pulp_write32(axi_m, 32'h6600193c, 32'h800003d4);
pulp_write32(axi_m, 32'h66001940, 32'h80000a64);
pulp_write32(axi_m, 32'h660000d8, 32'h00010000);
pulp_write32(axi_m, 32'h660000dc, 32'h00010001);
pulp_write32(axi_m, 32'h660000e0, 32'h00010002);
pulp_write32(axi_m, 32'h660000e4, 32'h00010003);
pulp_write32(axi_m, 32'h660000e8, 32'h00010004);
pulp_write32(axi_m, 32'h660000ec, 32'h00010005);
pulp_write32(axi_m, 32'h660000f0, 32'h00010006);
pulp_write32(axi_m, 32'h660000f4, 32'h00010007);
pulp_write32(axi_m, 32'h660000f8, 32'h00010008);
pulp_write32(axi_m, 32'h660000fc, 32'h00010009);
pulp_write32(axi_m, 32'h66000100, 32'h0001000a);
pulp_write32(axi_m, 32'h66000104, 32'h0001000b);
pulp_write32(axi_m, 32'h66000108, 32'h0001000c);
pulp_write32(axi_m, 32'h6600010c, 32'h0001000d);
pulp_write32(axi_m, 32'h66000110, 32'h0001000e);
pulp_write32(axi_m, 32'h66000114, 32'h0001000f);

pulp_write32(axi_m, 32'h66000118, 32'd2);
pulp_write32(axi_m, 32'h6600011c, 32'd2);
pulp_write32(axi_m, 32'h66000120, 32'h80001948);
pulp_write32(axi_m, 32'h66001948, 32'h800001a4);
pulp_write32(axi_m, 32'h6600194c, 32'h8000166c);
pulp_write32(axi_m, 32'h66000164, 32'h00020000);
pulp_write32(axi_m, 32'h66000168, 32'h00020001);
pulp_write32(axi_m, 32'h6600016c, 32'h00020002);
pulp_write32(axi_m, 32'h66000170, 32'h00020003);
pulp_write32(axi_m, 32'h66000174, 32'h00020004);
pulp_write32(axi_m, 32'h66000178, 32'h00020005);
pulp_write32(axi_m, 32'h6600017c, 32'h00020006);
pulp_write32(axi_m, 32'h66000180, 32'h00020007);
pulp_write32(axi_m, 32'h66000184, 32'h00020008);
pulp_write32(axi_m, 32'h66000188, 32'h00020009);
pulp_write32(axi_m, 32'h6600018c, 32'h0002000a);
pulp_write32(axi_m, 32'h66000190, 32'h0002000b);
pulp_write32(axi_m, 32'h66000194, 32'h0002000c);
pulp_write32(axi_m, 32'h66000198, 32'h0002000d);
pulp_write32(axi_m, 32'h6600019c, 32'h0002000e);
pulp_write32(axi_m, 32'h660001a0, 32'h0002000f);

pulp_write32(axi_m, 32'h660001a4, 32'd3);
pulp_write32(axi_m, 32'h660001a8, 32'd2);
pulp_write32(axi_m, 32'h660001ac, 32'h80001950);
pulp_write32(axi_m, 32'h66001950, 32'h80000230);
pulp_write32(axi_m, 32'h66001954, 32'h80000ec4);
pulp_write32(axi_m, 32'h660001f0, 32'h00030000);
pulp_write32(axi_m, 32'h660001f4, 32'h00030001);
pulp_write32(axi_m, 32'h660001f8, 32'h00030002);
pulp_write32(axi_m, 32'h660001fc, 32'h00030003);
pulp_write32(axi_m, 32'h66000200, 32'h00030004);
pulp_write32(axi_m, 32'h66000204, 32'h00030005);
pulp_write32(axi_m, 32'h66000208, 32'h00030006);
pulp_write32(axi_m, 32'h6600020c, 32'h00030007);
pulp_write32(axi_m, 32'h66000210, 32'h00030008);
pulp_write32(axi_m, 32'h66000214, 32'h00030009);
pulp_write32(axi_m, 32'h66000218, 32'h0003000a);
pulp_write32(axi_m, 32'h6600021c, 32'h0003000b);
pulp_write32(axi_m, 32'h66000220, 32'h0003000c);
pulp_write32(axi_m, 32'h66000224, 32'h0003000d);
pulp_write32(axi_m, 32'h66000228, 32'h0003000e);
pulp_write32(axi_m, 32'h6600022c, 32'h0003000f);

pulp_write32(axi_m, 32'h66000230, 32'd4);
pulp_write32(axi_m, 32'h66000234, 32'd2);
pulp_write32(axi_m, 32'h66000238, 32'h80001958);
pulp_write32(axi_m, 32'h66001958, 32'h800002bc);
pulp_write32(axi_m, 32'h6600195c, 32'h8000120c);
pulp_write32(axi_m, 32'h6600027c, 32'h00040000);
pulp_write32(axi_m, 32'h66000280, 32'h00040001);
pulp_write32(axi_m, 32'h66000284, 32'h00040002);
pulp_write32(axi_m, 32'h66000288, 32'h00040003);
pulp_write32(axi_m, 32'h6600028c, 32'h00040004);
pulp_write32(axi_m, 32'h66000290, 32'h00040005);
pulp_write32(axi_m, 32'h66000294, 32'h00040006);
pulp_write32(axi_m, 32'h66000298, 32'h00040007);
pulp_write32(axi_m, 32'h6600029c, 32'h00040008);
pulp_write32(axi_m, 32'h660002a0, 32'h00040009);
pulp_write32(axi_m, 32'h660002a4, 32'h0004000a);
pulp_write32(axi_m, 32'h660002a8, 32'h0004000b);
pulp_write32(axi_m, 32'h660002ac, 32'h0004000c);
pulp_write32(axi_m, 32'h660002b0, 32'h0004000d);
pulp_write32(axi_m, 32'h660002b4, 32'h0004000e);
pulp_write32(axi_m, 32'h660002b8, 32'h0004000f);

pulp_write32(axi_m, 32'h660002bc, 32'd5);
pulp_write32(axi_m, 32'h660002c0, 32'd2);
pulp_write32(axi_m, 32'h660002c4, 32'h80001960);
pulp_write32(axi_m, 32'h66001960, 32'h80000348);
pulp_write32(axi_m, 32'h66001964, 32'h8000189c);
pulp_write32(axi_m, 32'h66000308, 32'h00050000);
pulp_write32(axi_m, 32'h6600030c, 32'h00050001);
pulp_write32(axi_m, 32'h66000310, 32'h00050002);
pulp_write32(axi_m, 32'h66000314, 32'h00050003);
pulp_write32(axi_m, 32'h66000318, 32'h00050004);
pulp_write32(axi_m, 32'h6600031c, 32'h00050005);
pulp_write32(axi_m, 32'h66000320, 32'h00050006);
pulp_write32(axi_m, 32'h66000324, 32'h00050007);
pulp_write32(axi_m, 32'h66000328, 32'h00050008);
pulp_write32(axi_m, 32'h6600032c, 32'h00050009);
pulp_write32(axi_m, 32'h66000330, 32'h0005000a);
pulp_write32(axi_m, 32'h66000334, 32'h0005000b);
pulp_write32(axi_m, 32'h66000338, 32'h0005000c);
pulp_write32(axi_m, 32'h6600033c, 32'h0005000d);
pulp_write32(axi_m, 32'h66000340, 32'h0005000e);
pulp_write32(axi_m, 32'h66000344, 32'h0005000f);

pulp_write32(axi_m, 32'h66000348, 32'd6);
pulp_write32(axi_m, 32'h6600034c, 32'd2);
pulp_write32(axi_m, 32'h66000350, 32'h80001968);
pulp_write32(axi_m, 32'h66001968, 32'h800004ec);
pulp_write32(axi_m, 32'h6600196c, 32'h80000fdc);
pulp_write32(axi_m, 32'h66000394, 32'h00060000);
pulp_write32(axi_m, 32'h66000398, 32'h00060001);
pulp_write32(axi_m, 32'h6600039c, 32'h00060002);
pulp_write32(axi_m, 32'h660003a0, 32'h00060003);
pulp_write32(axi_m, 32'h660003a4, 32'h00060004);
pulp_write32(axi_m, 32'h660003a8, 32'h00060005);
pulp_write32(axi_m, 32'h660003ac, 32'h00060006);
pulp_write32(axi_m, 32'h660003b0, 32'h00060007);
pulp_write32(axi_m, 32'h660003b4, 32'h00060008);
pulp_write32(axi_m, 32'h660003b8, 32'h00060009);
pulp_write32(axi_m, 32'h660003bc, 32'h0006000a);
pulp_write32(axi_m, 32'h660003c0, 32'h0006000b);
pulp_write32(axi_m, 32'h660003c4, 32'h0006000c);
pulp_write32(axi_m, 32'h660003c8, 32'h0006000d);
pulp_write32(axi_m, 32'h660003cc, 32'h0006000e);
pulp_write32(axi_m, 32'h660003d0, 32'h0006000f);

pulp_write32(axi_m, 32'h660003d4, 32'd7);
pulp_write32(axi_m, 32'h660003d8, 32'd2);
pulp_write32(axi_m, 32'h660003dc, 32'h80001970);
pulp_write32(axi_m, 32'h66001970, 32'h80000460);
pulp_write32(axi_m, 32'h66001974, 32'h80000b7c);
pulp_write32(axi_m, 32'h66000420, 32'h00070000);
pulp_write32(axi_m, 32'h66000424, 32'h00070001);
pulp_write32(axi_m, 32'h66000428, 32'h00070002);
pulp_write32(axi_m, 32'h6600042c, 32'h00070003);
pulp_write32(axi_m, 32'h66000430, 32'h00070004);
pulp_write32(axi_m, 32'h66000434, 32'h00070005);
pulp_write32(axi_m, 32'h66000438, 32'h00070006);
pulp_write32(axi_m, 32'h6600043c, 32'h00070007);
pulp_write32(axi_m, 32'h66000440, 32'h00070008);
pulp_write32(axi_m, 32'h66000444, 32'h00070009);
pulp_write32(axi_m, 32'h66000448, 32'h0007000a);
pulp_write32(axi_m, 32'h6600044c, 32'h0007000b);
pulp_write32(axi_m, 32'h66000450, 32'h0007000c);
pulp_write32(axi_m, 32'h66000454, 32'h0007000d);
pulp_write32(axi_m, 32'h66000458, 32'h0007000e);
pulp_write32(axi_m, 32'h6600045c, 32'h0007000f);

pulp_write32(axi_m, 32'h66000460, 32'd8);
pulp_write32(axi_m, 32'h66000464, 32'd2);
pulp_write32(axi_m, 32'h66000468, 32'h80001978);
pulp_write32(axi_m, 32'h66001978, 32'h800004ec);
pulp_write32(axi_m, 32'h6600197c, 32'h80000c08);
pulp_write32(axi_m, 32'h660004ac, 32'h00080000);
pulp_write32(axi_m, 32'h660004b0, 32'h00080001);
pulp_write32(axi_m, 32'h660004b4, 32'h00080002);
pulp_write32(axi_m, 32'h660004b8, 32'h00080003);
pulp_write32(axi_m, 32'h660004bc, 32'h00080004);
pulp_write32(axi_m, 32'h660004c0, 32'h00080005);
pulp_write32(axi_m, 32'h660004c4, 32'h00080006);
pulp_write32(axi_m, 32'h660004c8, 32'h00080007);
pulp_write32(axi_m, 32'h660004cc, 32'h00080008);
pulp_write32(axi_m, 32'h660004d0, 32'h00080009);
pulp_write32(axi_m, 32'h660004d4, 32'h0008000a);
pulp_write32(axi_m, 32'h660004d8, 32'h0008000b);
pulp_write32(axi_m, 32'h660004dc, 32'h0008000c);
pulp_write32(axi_m, 32'h660004e0, 32'h0008000d);
pulp_write32(axi_m, 32'h660004e4, 32'h0008000e);
pulp_write32(axi_m, 32'h660004e8, 32'h0008000f);

pulp_write32(axi_m, 32'h660004ec, 32'd9);
pulp_write32(axi_m, 32'h660004f0, 32'd1);
pulp_write32(axi_m, 32'h660004f4, 32'h80001980);
pulp_write32(axi_m, 32'h66001980, 32'h80000d20);
pulp_write32(axi_m, 32'h66000538, 32'h00090000);
pulp_write32(axi_m, 32'h6600053c, 32'h00090001);
pulp_write32(axi_m, 32'h66000540, 32'h00090002);
pulp_write32(axi_m, 32'h66000544, 32'h00090003);
pulp_write32(axi_m, 32'h66000548, 32'h00090004);
pulp_write32(axi_m, 32'h6600054c, 32'h00090005);
pulp_write32(axi_m, 32'h66000550, 32'h00090006);
pulp_write32(axi_m, 32'h66000554, 32'h00090007);
pulp_write32(axi_m, 32'h66000558, 32'h00090008);
pulp_write32(axi_m, 32'h6600055c, 32'h00090009);
pulp_write32(axi_m, 32'h66000560, 32'h0009000a);
pulp_write32(axi_m, 32'h66000564, 32'h0009000b);
pulp_write32(axi_m, 32'h66000568, 32'h0009000c);
pulp_write32(axi_m, 32'h6600056c, 32'h0009000d);
pulp_write32(axi_m, 32'h66000570, 32'h0009000e);
pulp_write32(axi_m, 32'h66000574, 32'h0009000f);

pulp_write32(axi_m, 32'h66000578, 32'd10);
pulp_write32(axi_m, 32'h6600057c, 32'd2);
pulp_write32(axi_m, 32'h66000580, 32'h80001988);
pulp_write32(axi_m, 32'h66001988, 32'h8000071c);
pulp_write32(axi_m, 32'h6600198c, 32'h800007a8);
pulp_write32(axi_m, 32'h660005c4, 32'h000a0000);
pulp_write32(axi_m, 32'h660005c8, 32'h000a0001);
pulp_write32(axi_m, 32'h660005cc, 32'h000a0002);
pulp_write32(axi_m, 32'h660005d0, 32'h000a0003);
pulp_write32(axi_m, 32'h660005d4, 32'h000a0004);
pulp_write32(axi_m, 32'h660005d8, 32'h000a0005);
pulp_write32(axi_m, 32'h660005dc, 32'h000a0006);
pulp_write32(axi_m, 32'h660005e0, 32'h000a0007);
pulp_write32(axi_m, 32'h660005e4, 32'h000a0008);
pulp_write32(axi_m, 32'h660005e8, 32'h000a0009);
pulp_write32(axi_m, 32'h660005ec, 32'h000a000a);
pulp_write32(axi_m, 32'h660005f0, 32'h000a000b);
pulp_write32(axi_m, 32'h660005f4, 32'h000a000c);
pulp_write32(axi_m, 32'h660005f8, 32'h000a000d);
pulp_write32(axi_m, 32'h660005fc, 32'h000a000e);
pulp_write32(axi_m, 32'h66000600, 32'h000a000f);

pulp_write32(axi_m, 32'h66000604, 32'd11);
pulp_write32(axi_m, 32'h66000608, 32'd2);
pulp_write32(axi_m, 32'h6600060c, 32'h80001990);
pulp_write32(axi_m, 32'h66001990, 32'h80000e38);
pulp_write32(axi_m, 32'h66001994, 32'h80000f50);
pulp_write32(axi_m, 32'h66000650, 32'h000b0000);
pulp_write32(axi_m, 32'h66000654, 32'h000b0001);
pulp_write32(axi_m, 32'h66000658, 32'h000b0002);
pulp_write32(axi_m, 32'h6600065c, 32'h000b0003);
pulp_write32(axi_m, 32'h66000660, 32'h000b0004);
pulp_write32(axi_m, 32'h66000664, 32'h000b0005);
pulp_write32(axi_m, 32'h66000668, 32'h000b0006);
pulp_write32(axi_m, 32'h6600066c, 32'h000b0007);
pulp_write32(axi_m, 32'h66000670, 32'h000b0008);
pulp_write32(axi_m, 32'h66000674, 32'h000b0009);
pulp_write32(axi_m, 32'h66000678, 32'h000b000a);
pulp_write32(axi_m, 32'h6600067c, 32'h000b000b);
pulp_write32(axi_m, 32'h66000680, 32'h000b000c);
pulp_write32(axi_m, 32'h66000684, 32'h000b000d);
pulp_write32(axi_m, 32'h66000688, 32'h000b000e);
pulp_write32(axi_m, 32'h6600068c, 32'h000b000f);

pulp_write32(axi_m, 32'h66000690, 32'd12);
pulp_write32(axi_m, 32'h66000694, 32'd2);
pulp_write32(axi_m, 32'h66000698, 32'h80001998);
pulp_write32(axi_m, 32'h66001998, 32'h80001068);
pulp_write32(axi_m, 32'h6600199c, 32'h800010f4);
pulp_write32(axi_m, 32'h660006dc, 32'h000c0000);
pulp_write32(axi_m, 32'h660006e0, 32'h000c0001);
pulp_write32(axi_m, 32'h660006e4, 32'h000c0002);
pulp_write32(axi_m, 32'h660006e8, 32'h000c0003);
pulp_write32(axi_m, 32'h660006ec, 32'h000c0004);
pulp_write32(axi_m, 32'h660006f0, 32'h000c0005);
pulp_write32(axi_m, 32'h660006f4, 32'h000c0006);
pulp_write32(axi_m, 32'h660006f8, 32'h000c0007);
pulp_write32(axi_m, 32'h660006fc, 32'h000c0008);
pulp_write32(axi_m, 32'h66000700, 32'h000c0009);
pulp_write32(axi_m, 32'h66000704, 32'h000c000a);
pulp_write32(axi_m, 32'h66000708, 32'h000c000b);
pulp_write32(axi_m, 32'h6600070c, 32'h000c000c);
pulp_write32(axi_m, 32'h66000710, 32'h000c000d);
pulp_write32(axi_m, 32'h66000714, 32'h000c000e);
pulp_write32(axi_m, 32'h66000718, 32'h000c000f);

pulp_write32(axi_m, 32'h6600071c, 32'd13);
pulp_write32(axi_m, 32'h66000720, 32'd2);
pulp_write32(axi_m, 32'h66000724, 32'h800019a0);
pulp_write32(axi_m, 32'h660019a0, 32'h80000834);
pulp_write32(axi_m, 32'h660019a4, 32'h80000b7c);
pulp_write32(axi_m, 32'h66000768, 32'h000d0000);
pulp_write32(axi_m, 32'h6600076c, 32'h000d0001);
pulp_write32(axi_m, 32'h66000770, 32'h000d0002);
pulp_write32(axi_m, 32'h66000774, 32'h000d0003);
pulp_write32(axi_m, 32'h66000778, 32'h000d0004);
pulp_write32(axi_m, 32'h6600077c, 32'h000d0005);
pulp_write32(axi_m, 32'h66000780, 32'h000d0006);
pulp_write32(axi_m, 32'h66000784, 32'h000d0007);
pulp_write32(axi_m, 32'h66000788, 32'h000d0008);
pulp_write32(axi_m, 32'h6600078c, 32'h000d0009);
pulp_write32(axi_m, 32'h66000790, 32'h000d000a);
pulp_write32(axi_m, 32'h66000794, 32'h000d000b);
pulp_write32(axi_m, 32'h66000798, 32'h000d000c);
pulp_write32(axi_m, 32'h6600079c, 32'h000d000d);
pulp_write32(axi_m, 32'h660007a0, 32'h000d000e);
pulp_write32(axi_m, 32'h660007a4, 32'h000d000f);

pulp_write32(axi_m, 32'h660007a8, 32'd14);
pulp_write32(axi_m, 32'h660007ac, 32'd2);
pulp_write32(axi_m, 32'h660007b0, 32'h800019a8);
pulp_write32(axi_m, 32'h660019a8, 32'h80000834);
pulp_write32(axi_m, 32'h660019ac, 32'h800009d8);
pulp_write32(axi_m, 32'h660007f4, 32'h000e0000);
pulp_write32(axi_m, 32'h660007f8, 32'h000e0001);
pulp_write32(axi_m, 32'h660007fc, 32'h000e0002);
pulp_write32(axi_m, 32'h66000800, 32'h000e0003);
pulp_write32(axi_m, 32'h66000804, 32'h000e0004);
pulp_write32(axi_m, 32'h66000808, 32'h000e0005);
pulp_write32(axi_m, 32'h6600080c, 32'h000e0006);
pulp_write32(axi_m, 32'h66000810, 32'h000e0007);
pulp_write32(axi_m, 32'h66000814, 32'h000e0008);
pulp_write32(axi_m, 32'h66000818, 32'h000e0009);
pulp_write32(axi_m, 32'h6600081c, 32'h000e000a);
pulp_write32(axi_m, 32'h66000820, 32'h000e000b);
pulp_write32(axi_m, 32'h66000824, 32'h000e000c);
pulp_write32(axi_m, 32'h66000828, 32'h000e000d);
pulp_write32(axi_m, 32'h6600082c, 32'h000e000e);
pulp_write32(axi_m, 32'h66000830, 32'h000e000f);

pulp_write32(axi_m, 32'h66000834, 32'd15);
pulp_write32(axi_m, 32'h66000838, 32'd1);
pulp_write32(axi_m, 32'h6600083c, 32'h800019b0);
pulp_write32(axi_m, 32'h660019b0, 32'h800008c0);
pulp_write32(axi_m, 32'h66000880, 32'h000f0000);
pulp_write32(axi_m, 32'h66000884, 32'h000f0001);
pulp_write32(axi_m, 32'h66000888, 32'h000f0002);
pulp_write32(axi_m, 32'h6600088c, 32'h000f0003);
pulp_write32(axi_m, 32'h66000890, 32'h000f0004);
pulp_write32(axi_m, 32'h66000894, 32'h000f0005);
pulp_write32(axi_m, 32'h66000898, 32'h000f0006);
pulp_write32(axi_m, 32'h6600089c, 32'h000f0007);
pulp_write32(axi_m, 32'h660008a0, 32'h000f0008);
pulp_write32(axi_m, 32'h660008a4, 32'h000f0009);
pulp_write32(axi_m, 32'h660008a8, 32'h000f000a);
pulp_write32(axi_m, 32'h660008ac, 32'h000f000b);
pulp_write32(axi_m, 32'h660008b0, 32'h000f000c);
pulp_write32(axi_m, 32'h660008b4, 32'h000f000d);
pulp_write32(axi_m, 32'h660008b8, 32'h000f000e);
pulp_write32(axi_m, 32'h660008bc, 32'h000f000f);

pulp_write32(axi_m, 32'h660008c0, 32'd16);
pulp_write32(axi_m, 32'h660008c4, 32'd2);
pulp_write32(axi_m, 32'h660008c8, 32'h800019b8);
pulp_write32(axi_m, 32'h660019b8, 32'h8000094c);
pulp_write32(axi_m, 32'h660019bc, 32'h80000af0);
pulp_write32(axi_m, 32'h6600090c, 32'h00100000);
pulp_write32(axi_m, 32'h66000910, 32'h00100001);
pulp_write32(axi_m, 32'h66000914, 32'h00100002);
pulp_write32(axi_m, 32'h66000918, 32'h00100003);
pulp_write32(axi_m, 32'h6600091c, 32'h00100004);
pulp_write32(axi_m, 32'h66000920, 32'h00100005);
pulp_write32(axi_m, 32'h66000924, 32'h00100006);
pulp_write32(axi_m, 32'h66000928, 32'h00100007);
pulp_write32(axi_m, 32'h6600092c, 32'h00100008);
pulp_write32(axi_m, 32'h66000930, 32'h00100009);
pulp_write32(axi_m, 32'h66000934, 32'h0010000a);
pulp_write32(axi_m, 32'h66000938, 32'h0010000b);
pulp_write32(axi_m, 32'h6600093c, 32'h0010000c);
pulp_write32(axi_m, 32'h66000940, 32'h0010000d);
pulp_write32(axi_m, 32'h66000944, 32'h0010000e);
pulp_write32(axi_m, 32'h66000948, 32'h0010000f);

pulp_write32(axi_m, 32'h6600094c, 32'd17);
pulp_write32(axi_m, 32'h66000950, 32'd2);
pulp_write32(axi_m, 32'h66000954, 32'h800019c0);
pulp_write32(axi_m, 32'h660019c0, 32'h800009d8);
pulp_write32(axi_m, 32'h660019c4, 32'h80000c94);
pulp_write32(axi_m, 32'h66000998, 32'h00110000);
pulp_write32(axi_m, 32'h6600099c, 32'h00110001);
pulp_write32(axi_m, 32'h660009a0, 32'h00110002);
pulp_write32(axi_m, 32'h660009a4, 32'h00110003);
pulp_write32(axi_m, 32'h660009a8, 32'h00110004);
pulp_write32(axi_m, 32'h660009ac, 32'h00110005);
pulp_write32(axi_m, 32'h660009b0, 32'h00110006);
pulp_write32(axi_m, 32'h660009b4, 32'h00110007);
pulp_write32(axi_m, 32'h660009b8, 32'h00110008);
pulp_write32(axi_m, 32'h660009bc, 32'h00110009);
pulp_write32(axi_m, 32'h660009c0, 32'h0011000a);
pulp_write32(axi_m, 32'h660009c4, 32'h0011000b);
pulp_write32(axi_m, 32'h660009c8, 32'h0011000c);
pulp_write32(axi_m, 32'h660009cc, 32'h0011000d);
pulp_write32(axi_m, 32'h660009d0, 32'h0011000e);
pulp_write32(axi_m, 32'h660009d4, 32'h0011000f);

pulp_write32(axi_m, 32'h660009d8, 32'd18);
pulp_write32(axi_m, 32'h660009dc, 32'd1);
pulp_write32(axi_m, 32'h660009e0, 32'h800019c8);
pulp_write32(axi_m, 32'h660019c8, 32'h80000d20);
pulp_write32(axi_m, 32'h66000a24, 32'h00120000);
pulp_write32(axi_m, 32'h66000a28, 32'h00120001);
pulp_write32(axi_m, 32'h66000a2c, 32'h00120002);
pulp_write32(axi_m, 32'h66000a30, 32'h00120003);
pulp_write32(axi_m, 32'h66000a34, 32'h00120004);
pulp_write32(axi_m, 32'h66000a38, 32'h00120005);
pulp_write32(axi_m, 32'h66000a3c, 32'h00120006);
pulp_write32(axi_m, 32'h66000a40, 32'h00120007);
pulp_write32(axi_m, 32'h66000a44, 32'h00120008);
pulp_write32(axi_m, 32'h66000a48, 32'h00120009);
pulp_write32(axi_m, 32'h66000a4c, 32'h0012000a);
pulp_write32(axi_m, 32'h66000a50, 32'h0012000b);
pulp_write32(axi_m, 32'h66000a54, 32'h0012000c);
pulp_write32(axi_m, 32'h66000a58, 32'h0012000d);
pulp_write32(axi_m, 32'h66000a5c, 32'h0012000e);
pulp_write32(axi_m, 32'h66000a60, 32'h0012000f);

pulp_write32(axi_m, 32'h66000a64, 32'd19);
pulp_write32(axi_m, 32'h66000a68, 32'd2);
pulp_write32(axi_m, 32'h66000a6c, 32'h800019d0);
pulp_write32(axi_m, 32'h660019d0, 32'h80000dac);
pulp_write32(axi_m, 32'h660019d4, 32'h800015e0);
pulp_write32(axi_m, 32'h66000ab0, 32'h00130000);
pulp_write32(axi_m, 32'h66000ab4, 32'h00130001);
pulp_write32(axi_m, 32'h66000ab8, 32'h00130002);
pulp_write32(axi_m, 32'h66000abc, 32'h00130003);
pulp_write32(axi_m, 32'h66000ac0, 32'h00130004);
pulp_write32(axi_m, 32'h66000ac4, 32'h00130005);
pulp_write32(axi_m, 32'h66000ac8, 32'h00130006);
pulp_write32(axi_m, 32'h66000acc, 32'h00130007);
pulp_write32(axi_m, 32'h66000ad0, 32'h00130008);
pulp_write32(axi_m, 32'h66000ad4, 32'h00130009);
pulp_write32(axi_m, 32'h66000ad8, 32'h0013000a);
pulp_write32(axi_m, 32'h66000adc, 32'h0013000b);
pulp_write32(axi_m, 32'h66000ae0, 32'h0013000c);
pulp_write32(axi_m, 32'h66000ae4, 32'h0013000d);
pulp_write32(axi_m, 32'h66000ae8, 32'h0013000e);
pulp_write32(axi_m, 32'h66000aec, 32'h0013000f);

pulp_write32(axi_m, 32'h66000af0, 32'd20);
pulp_write32(axi_m, 32'h66000af4, 32'd2);
pulp_write32(axi_m, 32'h66000af8, 32'h800019d8);
pulp_write32(axi_m, 32'h660019d8, 32'h80000b7c);
pulp_write32(axi_m, 32'h660019dc, 32'h80000c08);
pulp_write32(axi_m, 32'h66000b3c, 32'h00140000);
pulp_write32(axi_m, 32'h66000b40, 32'h00140001);
pulp_write32(axi_m, 32'h66000b44, 32'h00140002);
pulp_write32(axi_m, 32'h66000b48, 32'h00140003);
pulp_write32(axi_m, 32'h66000b4c, 32'h00140004);
pulp_write32(axi_m, 32'h66000b50, 32'h00140005);
pulp_write32(axi_m, 32'h66000b54, 32'h00140006);
pulp_write32(axi_m, 32'h66000b58, 32'h00140007);
pulp_write32(axi_m, 32'h66000b5c, 32'h00140008);
pulp_write32(axi_m, 32'h66000b60, 32'h00140009);
pulp_write32(axi_m, 32'h66000b64, 32'h0014000a);
pulp_write32(axi_m, 32'h66000b68, 32'h0014000b);
pulp_write32(axi_m, 32'h66000b6c, 32'h0014000c);
pulp_write32(axi_m, 32'h66000b70, 32'h0014000d);
pulp_write32(axi_m, 32'h66000b74, 32'h0014000e);
pulp_write32(axi_m, 32'h66000b78, 32'h0014000f);

pulp_write32(axi_m, 32'h66000b7c, 32'd21);
pulp_write32(axi_m, 32'h66000b80, 32'd0);
pulp_write32(axi_m, 32'h66000bc8, 32'h00150000);
pulp_write32(axi_m, 32'h66000bcc, 32'h00150001);
pulp_write32(axi_m, 32'h66000bd0, 32'h00150002);
pulp_write32(axi_m, 32'h66000bd4, 32'h00150003);
pulp_write32(axi_m, 32'h66000bd8, 32'h00150004);
pulp_write32(axi_m, 32'h66000bdc, 32'h00150005);
pulp_write32(axi_m, 32'h66000be0, 32'h00150006);
pulp_write32(axi_m, 32'h66000be4, 32'h00150007);
pulp_write32(axi_m, 32'h66000be8, 32'h00150008);
pulp_write32(axi_m, 32'h66000bec, 32'h00150009);
pulp_write32(axi_m, 32'h66000bf0, 32'h0015000a);
pulp_write32(axi_m, 32'h66000bf4, 32'h0015000b);
pulp_write32(axi_m, 32'h66000bf8, 32'h0015000c);
pulp_write32(axi_m, 32'h66000bfc, 32'h0015000d);
pulp_write32(axi_m, 32'h66000c00, 32'h0015000e);
pulp_write32(axi_m, 32'h66000c04, 32'h0015000f);

pulp_write32(axi_m, 32'h66000c08, 32'd22);
pulp_write32(axi_m, 32'h66000c0c, 32'd1);
pulp_write32(axi_m, 32'h66000c10, 32'h800019e0);
pulp_write32(axi_m, 32'h660019e0, 32'h80000c94);
pulp_write32(axi_m, 32'h66000c54, 32'h00160000);
pulp_write32(axi_m, 32'h66000c58, 32'h00160001);
pulp_write32(axi_m, 32'h66000c5c, 32'h00160002);
pulp_write32(axi_m, 32'h66000c60, 32'h00160003);
pulp_write32(axi_m, 32'h66000c64, 32'h00160004);
pulp_write32(axi_m, 32'h66000c68, 32'h00160005);
pulp_write32(axi_m, 32'h66000c6c, 32'h00160006);
pulp_write32(axi_m, 32'h66000c70, 32'h00160007);
pulp_write32(axi_m, 32'h66000c74, 32'h00160008);
pulp_write32(axi_m, 32'h66000c78, 32'h00160009);
pulp_write32(axi_m, 32'h66000c7c, 32'h0016000a);
pulp_write32(axi_m, 32'h66000c80, 32'h0016000b);
pulp_write32(axi_m, 32'h66000c84, 32'h0016000c);
pulp_write32(axi_m, 32'h66000c88, 32'h0016000d);
pulp_write32(axi_m, 32'h66000c8c, 32'h0016000e);
pulp_write32(axi_m, 32'h66000c90, 32'h0016000f);

pulp_write32(axi_m, 32'h66000c94, 32'd23);
pulp_write32(axi_m, 32'h66000c98, 32'd1);
pulp_write32(axi_m, 32'h66000c9c, 32'h800019e8);
pulp_write32(axi_m, 32'h660019e8, 32'h80000d20);
pulp_write32(axi_m, 32'h66000ce0, 32'h00170000);
pulp_write32(axi_m, 32'h66000ce4, 32'h00170001);
pulp_write32(axi_m, 32'h66000ce8, 32'h00170002);
pulp_write32(axi_m, 32'h66000cec, 32'h00170003);
pulp_write32(axi_m, 32'h66000cf0, 32'h00170004);
pulp_write32(axi_m, 32'h66000cf4, 32'h00170005);
pulp_write32(axi_m, 32'h66000cf8, 32'h00170006);
pulp_write32(axi_m, 32'h66000cfc, 32'h00170007);
pulp_write32(axi_m, 32'h66000d00, 32'h00170008);
pulp_write32(axi_m, 32'h66000d04, 32'h00170009);
pulp_write32(axi_m, 32'h66000d08, 32'h0017000a);
pulp_write32(axi_m, 32'h66000d0c, 32'h0017000b);
pulp_write32(axi_m, 32'h66000d10, 32'h0017000c);
pulp_write32(axi_m, 32'h66000d14, 32'h0017000d);
pulp_write32(axi_m, 32'h66000d18, 32'h0017000e);
pulp_write32(axi_m, 32'h66000d1c, 32'h0017000f);

pulp_write32(axi_m, 32'h66000d20, 32'd24);
pulp_write32(axi_m, 32'h66000d24, 32'd0);
pulp_write32(axi_m, 32'h66000d6c, 32'h00180000);
pulp_write32(axi_m, 32'h66000d70, 32'h00180001);
pulp_write32(axi_m, 32'h66000d74, 32'h00180002);
pulp_write32(axi_m, 32'h66000d78, 32'h00180003);
pulp_write32(axi_m, 32'h66000d7c, 32'h00180004);
pulp_write32(axi_m, 32'h66000d80, 32'h00180005);
pulp_write32(axi_m, 32'h66000d84, 32'h00180006);
pulp_write32(axi_m, 32'h66000d88, 32'h00180007);
pulp_write32(axi_m, 32'h66000d8c, 32'h00180008);
pulp_write32(axi_m, 32'h66000d90, 32'h00180009);
pulp_write32(axi_m, 32'h66000d94, 32'h0018000a);
pulp_write32(axi_m, 32'h66000d98, 32'h0018000b);
pulp_write32(axi_m, 32'h66000d9c, 32'h0018000c);
pulp_write32(axi_m, 32'h66000da0, 32'h0018000d);
pulp_write32(axi_m, 32'h66000da4, 32'h0018000e);
pulp_write32(axi_m, 32'h66000da8, 32'h0018000f);

pulp_write32(axi_m, 32'h66000dac, 32'd25);
pulp_write32(axi_m, 32'h66000db0, 32'd2);
pulp_write32(axi_m, 32'h66000db4, 32'h800019f0);
pulp_write32(axi_m, 32'h660019f0, 32'h80000e38);
pulp_write32(axi_m, 32'h660019f4, 32'h800014c8);
pulp_write32(axi_m, 32'h66000df8, 32'h00190000);
pulp_write32(axi_m, 32'h66000dfc, 32'h00190001);
pulp_write32(axi_m, 32'h66000e00, 32'h00190002);
pulp_write32(axi_m, 32'h66000e04, 32'h00190003);
pulp_write32(axi_m, 32'h66000e08, 32'h00190004);
pulp_write32(axi_m, 32'h66000e0c, 32'h00190005);
pulp_write32(axi_m, 32'h66000e10, 32'h00190006);
pulp_write32(axi_m, 32'h66000e14, 32'h00190007);
pulp_write32(axi_m, 32'h66000e18, 32'h00190008);
pulp_write32(axi_m, 32'h66000e1c, 32'h00190009);
pulp_write32(axi_m, 32'h66000e20, 32'h0019000a);
pulp_write32(axi_m, 32'h66000e24, 32'h0019000b);
pulp_write32(axi_m, 32'h66000e28, 32'h0019000c);
pulp_write32(axi_m, 32'h66000e2c, 32'h0019000d);
pulp_write32(axi_m, 32'h66000e30, 32'h0019000e);
pulp_write32(axi_m, 32'h66000e34, 32'h0019000f);

pulp_write32(axi_m, 32'h66000e38, 32'd26);
pulp_write32(axi_m, 32'h66000e3c, 32'd1);
pulp_write32(axi_m, 32'h66000e40, 32'h800019f8);
pulp_write32(axi_m, 32'h660019f8, 32'h80001298);
pulp_write32(axi_m, 32'h66000e84, 32'h001a0000);
pulp_write32(axi_m, 32'h66000e88, 32'h001a0001);
pulp_write32(axi_m, 32'h66000e8c, 32'h001a0002);
pulp_write32(axi_m, 32'h66000e90, 32'h001a0003);
pulp_write32(axi_m, 32'h66000e94, 32'h001a0004);
pulp_write32(axi_m, 32'h66000e98, 32'h001a0005);
pulp_write32(axi_m, 32'h66000e9c, 32'h001a0006);
pulp_write32(axi_m, 32'h66000ea0, 32'h001a0007);
pulp_write32(axi_m, 32'h66000ea4, 32'h001a0008);
pulp_write32(axi_m, 32'h66000ea8, 32'h001a0009);
pulp_write32(axi_m, 32'h66000eac, 32'h001a000a);
pulp_write32(axi_m, 32'h66000eb0, 32'h001a000b);
pulp_write32(axi_m, 32'h66000eb4, 32'h001a000c);
pulp_write32(axi_m, 32'h66000eb8, 32'h001a000d);
pulp_write32(axi_m, 32'h66000ebc, 32'h001a000e);
pulp_write32(axi_m, 32'h66000ec0, 32'h001a000f);

pulp_write32(axi_m, 32'h66000ec4, 32'd27);
pulp_write32(axi_m, 32'h66000ec8, 32'd2);
pulp_write32(axi_m, 32'h66000ecc, 32'h80001a00);
pulp_write32(axi_m, 32'h66001a00, 32'h80000f50);
pulp_write32(axi_m, 32'h66001a04, 32'h80001554);
pulp_write32(axi_m, 32'h66000f10, 32'h001b0000);
pulp_write32(axi_m, 32'h66000f14, 32'h001b0001);
pulp_write32(axi_m, 32'h66000f18, 32'h001b0002);
pulp_write32(axi_m, 32'h66000f1c, 32'h001b0003);
pulp_write32(axi_m, 32'h66000f20, 32'h001b0004);
pulp_write32(axi_m, 32'h66000f24, 32'h001b0005);
pulp_write32(axi_m, 32'h66000f28, 32'h001b0006);
pulp_write32(axi_m, 32'h66000f2c, 32'h001b0007);
pulp_write32(axi_m, 32'h66000f30, 32'h001b0008);
pulp_write32(axi_m, 32'h66000f34, 32'h001b0009);
pulp_write32(axi_m, 32'h66000f38, 32'h001b000a);
pulp_write32(axi_m, 32'h66000f3c, 32'h001b000b);
pulp_write32(axi_m, 32'h66000f40, 32'h001b000c);
pulp_write32(axi_m, 32'h66000f44, 32'h001b000d);
pulp_write32(axi_m, 32'h66000f48, 32'h001b000e);
pulp_write32(axi_m, 32'h66000f4c, 32'h001b000f);

pulp_write32(axi_m, 32'h66000f50, 32'd28);
pulp_write32(axi_m, 32'h66000f54, 32'd1);
pulp_write32(axi_m, 32'h66000f58, 32'h80001a08);
pulp_write32(axi_m, 32'h66001a08, 32'h80001298);
pulp_write32(axi_m, 32'h66000f9c, 32'h001c0000);
pulp_write32(axi_m, 32'h66000fa0, 32'h001c0001);
pulp_write32(axi_m, 32'h66000fa4, 32'h001c0002);
pulp_write32(axi_m, 32'h66000fa8, 32'h001c0003);
pulp_write32(axi_m, 32'h66000fac, 32'h001c0004);
pulp_write32(axi_m, 32'h66000fb0, 32'h001c0005);
pulp_write32(axi_m, 32'h66000fb4, 32'h001c0006);
pulp_write32(axi_m, 32'h66000fb8, 32'h001c0007);
pulp_write32(axi_m, 32'h66000fbc, 32'h001c0008);
pulp_write32(axi_m, 32'h66000fc0, 32'h001c0009);
pulp_write32(axi_m, 32'h66000fc4, 32'h001c000a);
pulp_write32(axi_m, 32'h66000fc8, 32'h001c000b);
pulp_write32(axi_m, 32'h66000fcc, 32'h001c000c);
pulp_write32(axi_m, 32'h66000fd0, 32'h001c000d);
pulp_write32(axi_m, 32'h66000fd4, 32'h001c000e);
pulp_write32(axi_m, 32'h66000fd8, 32'h001c000f);

pulp_write32(axi_m, 32'h66000fdc, 32'd29);
pulp_write32(axi_m, 32'h66000fe0, 32'd2);
pulp_write32(axi_m, 32'h66000fe4, 32'h80001a10);
pulp_write32(axi_m, 32'h66001a10, 32'h80001068);
pulp_write32(axi_m, 32'h66001a14, 32'h80001810);
pulp_write32(axi_m, 32'h66001028, 32'h001d0000);
pulp_write32(axi_m, 32'h6600102c, 32'h001d0001);
pulp_write32(axi_m, 32'h66001030, 32'h001d0002);
pulp_write32(axi_m, 32'h66001034, 32'h001d0003);
pulp_write32(axi_m, 32'h66001038, 32'h001d0004);
pulp_write32(axi_m, 32'h6600103c, 32'h001d0005);
pulp_write32(axi_m, 32'h66001040, 32'h001d0006);
pulp_write32(axi_m, 32'h66001044, 32'h001d0007);
pulp_write32(axi_m, 32'h66001048, 32'h001d0008);
pulp_write32(axi_m, 32'h6600104c, 32'h001d0009);
pulp_write32(axi_m, 32'h66001050, 32'h001d000a);
pulp_write32(axi_m, 32'h66001054, 32'h001d000b);
pulp_write32(axi_m, 32'h66001058, 32'h001d000c);
pulp_write32(axi_m, 32'h6600105c, 32'h001d000d);
pulp_write32(axi_m, 32'h66001060, 32'h001d000e);
pulp_write32(axi_m, 32'h66001064, 32'h001d000f);

pulp_write32(axi_m, 32'h66001068, 32'd30);
pulp_write32(axi_m, 32'h6600106c, 32'd1);
pulp_write32(axi_m, 32'h66001070, 32'h80001a18);
pulp_write32(axi_m, 32'h66001a18, 32'h80001324);
pulp_write32(axi_m, 32'h660010b4, 32'h001e0000);
pulp_write32(axi_m, 32'h660010b8, 32'h001e0001);
pulp_write32(axi_m, 32'h660010bc, 32'h001e0002);
pulp_write32(axi_m, 32'h660010c0, 32'h001e0003);
pulp_write32(axi_m, 32'h660010c4, 32'h001e0004);
pulp_write32(axi_m, 32'h660010c8, 32'h001e0005);
pulp_write32(axi_m, 32'h660010cc, 32'h001e0006);
pulp_write32(axi_m, 32'h660010d0, 32'h001e0007);
pulp_write32(axi_m, 32'h660010d4, 32'h001e0008);
pulp_write32(axi_m, 32'h660010d8, 32'h001e0009);
pulp_write32(axi_m, 32'h660010dc, 32'h001e000a);
pulp_write32(axi_m, 32'h660010e0, 32'h001e000b);
pulp_write32(axi_m, 32'h660010e4, 32'h001e000c);
pulp_write32(axi_m, 32'h660010e8, 32'h001e000d);
pulp_write32(axi_m, 32'h660010ec, 32'h001e000e);
pulp_write32(axi_m, 32'h660010f0, 32'h001e000f);

pulp_write32(axi_m, 32'h660010f4, 32'd31);
pulp_write32(axi_m, 32'h660010f8, 32'd2);
pulp_write32(axi_m, 32'h660010fc, 32'h80001a20);
pulp_write32(axi_m, 32'h66001a20, 32'h80001180);
pulp_write32(axi_m, 32'h66001a24, 32'h80001324);
pulp_write32(axi_m, 32'h66001140, 32'h001f0000);
pulp_write32(axi_m, 32'h66001144, 32'h001f0001);
pulp_write32(axi_m, 32'h66001148, 32'h001f0002);
pulp_write32(axi_m, 32'h6600114c, 32'h001f0003);
pulp_write32(axi_m, 32'h66001150, 32'h001f0004);
pulp_write32(axi_m, 32'h66001154, 32'h001f0005);
pulp_write32(axi_m, 32'h66001158, 32'h001f0006);
pulp_write32(axi_m, 32'h6600115c, 32'h001f0007);
pulp_write32(axi_m, 32'h66001160, 32'h001f0008);
pulp_write32(axi_m, 32'h66001164, 32'h001f0009);
pulp_write32(axi_m, 32'h66001168, 32'h001f000a);
pulp_write32(axi_m, 32'h6600116c, 32'h001f000b);
pulp_write32(axi_m, 32'h66001170, 32'h001f000c);
pulp_write32(axi_m, 32'h66001174, 32'h001f000d);
pulp_write32(axi_m, 32'h66001178, 32'h001f000e);
pulp_write32(axi_m, 32'h6600117c, 32'h001f000f);

pulp_write32(axi_m, 32'h66001180, 32'd32);
pulp_write32(axi_m, 32'h66001184, 32'd2);
pulp_write32(axi_m, 32'h66001188, 32'h80001a28);
pulp_write32(axi_m, 32'h66001a28, 32'h8000120c);
pulp_write32(axi_m, 32'h66001a2c, 32'h800016f8);
pulp_write32(axi_m, 32'h660011cc, 32'h00200000);
pulp_write32(axi_m, 32'h660011d0, 32'h00200001);
pulp_write32(axi_m, 32'h660011d4, 32'h00200002);
pulp_write32(axi_m, 32'h660011d8, 32'h00200003);
pulp_write32(axi_m, 32'h660011dc, 32'h00200004);
pulp_write32(axi_m, 32'h660011e0, 32'h00200005);
pulp_write32(axi_m, 32'h660011e4, 32'h00200006);
pulp_write32(axi_m, 32'h660011e8, 32'h00200007);
pulp_write32(axi_m, 32'h660011ec, 32'h00200008);
pulp_write32(axi_m, 32'h660011f0, 32'h00200009);
pulp_write32(axi_m, 32'h660011f4, 32'h0020000a);
pulp_write32(axi_m, 32'h660011f8, 32'h0020000b);
pulp_write32(axi_m, 32'h660011fc, 32'h0020000c);
pulp_write32(axi_m, 32'h66001200, 32'h0020000d);
pulp_write32(axi_m, 32'h66001204, 32'h0020000e);
pulp_write32(axi_m, 32'h66001208, 32'h0020000f);

pulp_write32(axi_m, 32'h6600120c, 32'd33);
pulp_write32(axi_m, 32'h66001210, 32'd1);
pulp_write32(axi_m, 32'h66001214, 32'h80001a30);
pulp_write32(axi_m, 32'h66001a30, 32'h80001784);
pulp_write32(axi_m, 32'h66001258, 32'h00210000);
pulp_write32(axi_m, 32'h6600125c, 32'h00210001);
pulp_write32(axi_m, 32'h66001260, 32'h00210002);
pulp_write32(axi_m, 32'h66001264, 32'h00210003);
pulp_write32(axi_m, 32'h66001268, 32'h00210004);
pulp_write32(axi_m, 32'h6600126c, 32'h00210005);
pulp_write32(axi_m, 32'h66001270, 32'h00210006);
pulp_write32(axi_m, 32'h66001274, 32'h00210007);
pulp_write32(axi_m, 32'h66001278, 32'h00210008);
pulp_write32(axi_m, 32'h6600127c, 32'h00210009);
pulp_write32(axi_m, 32'h66001280, 32'h0021000a);
pulp_write32(axi_m, 32'h66001284, 32'h0021000b);
pulp_write32(axi_m, 32'h66001288, 32'h0021000c);
pulp_write32(axi_m, 32'h6600128c, 32'h0021000d);
pulp_write32(axi_m, 32'h66001290, 32'h0021000e);
pulp_write32(axi_m, 32'h66001294, 32'h0021000f);

pulp_write32(axi_m, 32'h66001298, 32'd34);
pulp_write32(axi_m, 32'h6600129c, 32'd1);
pulp_write32(axi_m, 32'h660012a0, 32'h80001a38);
pulp_write32(axi_m, 32'h66001a38, 32'h800013b0);
pulp_write32(axi_m, 32'h660012e4, 32'h00220000);
pulp_write32(axi_m, 32'h660012e8, 32'h00220001);
pulp_write32(axi_m, 32'h660012ec, 32'h00220002);
pulp_write32(axi_m, 32'h660012f0, 32'h00220003);
pulp_write32(axi_m, 32'h660012f4, 32'h00220004);
pulp_write32(axi_m, 32'h660012f8, 32'h00220005);
pulp_write32(axi_m, 32'h660012fc, 32'h00220006);
pulp_write32(axi_m, 32'h66001300, 32'h00220007);
pulp_write32(axi_m, 32'h66001304, 32'h00220008);
pulp_write32(axi_m, 32'h66001308, 32'h00220009);
pulp_write32(axi_m, 32'h6600130c, 32'h0022000a);
pulp_write32(axi_m, 32'h66001310, 32'h0022000b);
pulp_write32(axi_m, 32'h66001314, 32'h0022000c);
pulp_write32(axi_m, 32'h66001318, 32'h0022000d);
pulp_write32(axi_m, 32'h6600131c, 32'h0022000e);
pulp_write32(axi_m, 32'h66001320, 32'h0022000f);

pulp_write32(axi_m, 32'h66001324, 32'd35);
pulp_write32(axi_m, 32'h66001328, 32'd1);
pulp_write32(axi_m, 32'h6600132c, 32'h80001a40);
pulp_write32(axi_m, 32'h66001a40, 32'h8000143c);
pulp_write32(axi_m, 32'h66001370, 32'h00230000);
pulp_write32(axi_m, 32'h66001374, 32'h00230001);
pulp_write32(axi_m, 32'h66001378, 32'h00230002);
pulp_write32(axi_m, 32'h6600137c, 32'h00230003);
pulp_write32(axi_m, 32'h66001380, 32'h00230004);
pulp_write32(axi_m, 32'h66001384, 32'h00230005);
pulp_write32(axi_m, 32'h66001388, 32'h00230006);
pulp_write32(axi_m, 32'h6600138c, 32'h00230007);
pulp_write32(axi_m, 32'h66001390, 32'h00230008);
pulp_write32(axi_m, 32'h66001394, 32'h00230009);
pulp_write32(axi_m, 32'h66001398, 32'h0023000a);
pulp_write32(axi_m, 32'h6600139c, 32'h0023000b);
pulp_write32(axi_m, 32'h660013a0, 32'h0023000c);
pulp_write32(axi_m, 32'h660013a4, 32'h0023000d);
pulp_write32(axi_m, 32'h660013a8, 32'h0023000e);
pulp_write32(axi_m, 32'h660013ac, 32'h0023000f);

pulp_write32(axi_m, 32'h660013b0, 32'd36);
pulp_write32(axi_m, 32'h660013b4, 32'd2);
pulp_write32(axi_m, 32'h660013b8, 32'h80001a48);
pulp_write32(axi_m, 32'h66001a48, 32'h800014c8);
pulp_write32(axi_m, 32'h66001a4c, 32'h80001554);
pulp_write32(axi_m, 32'h660013fc, 32'h00240000);
pulp_write32(axi_m, 32'h66001400, 32'h00240001);
pulp_write32(axi_m, 32'h66001404, 32'h00240002);
pulp_write32(axi_m, 32'h66001408, 32'h00240003);
pulp_write32(axi_m, 32'h6600140c, 32'h00240004);
pulp_write32(axi_m, 32'h66001410, 32'h00240005);
pulp_write32(axi_m, 32'h66001414, 32'h00240006);
pulp_write32(axi_m, 32'h66001418, 32'h00240007);
pulp_write32(axi_m, 32'h6600141c, 32'h00240008);
pulp_write32(axi_m, 32'h66001420, 32'h00240009);
pulp_write32(axi_m, 32'h66001424, 32'h0024000a);
pulp_write32(axi_m, 32'h66001428, 32'h0024000b);
pulp_write32(axi_m, 32'h6600142c, 32'h0024000c);
pulp_write32(axi_m, 32'h66001430, 32'h0024000d);
pulp_write32(axi_m, 32'h66001434, 32'h0024000e);
pulp_write32(axi_m, 32'h66001438, 32'h0024000f);

pulp_write32(axi_m, 32'h6600143c, 32'd37);
pulp_write32(axi_m, 32'h66001440, 32'd2);
pulp_write32(axi_m, 32'h66001444, 32'h80001a50);
pulp_write32(axi_m, 32'h66001a50, 32'h800016f8);
pulp_write32(axi_m, 32'h66001a54, 32'h80001810);
pulp_write32(axi_m, 32'h66001488, 32'h00250000);
pulp_write32(axi_m, 32'h6600148c, 32'h00250001);
pulp_write32(axi_m, 32'h66001490, 32'h00250002);
pulp_write32(axi_m, 32'h66001494, 32'h00250003);
pulp_write32(axi_m, 32'h66001498, 32'h00250004);
pulp_write32(axi_m, 32'h6600149c, 32'h00250005);
pulp_write32(axi_m, 32'h660014a0, 32'h00250006);
pulp_write32(axi_m, 32'h660014a4, 32'h00250007);
pulp_write32(axi_m, 32'h660014a8, 32'h00250008);
pulp_write32(axi_m, 32'h660014ac, 32'h00250009);
pulp_write32(axi_m, 32'h660014b0, 32'h0025000a);
pulp_write32(axi_m, 32'h660014b4, 32'h0025000b);
pulp_write32(axi_m, 32'h660014b8, 32'h0025000c);
pulp_write32(axi_m, 32'h660014bc, 32'h0025000d);
pulp_write32(axi_m, 32'h660014c0, 32'h0025000e);
pulp_write32(axi_m, 32'h660014c4, 32'h0025000f);

pulp_write32(axi_m, 32'h660014c8, 32'd38);
pulp_write32(axi_m, 32'h660014cc, 32'd1);
pulp_write32(axi_m, 32'h660014d0, 32'h80001a58);
pulp_write32(axi_m, 32'h66001a58, 32'h800015e0);
pulp_write32(axi_m, 32'h66001514, 32'h00260000);
pulp_write32(axi_m, 32'h66001518, 32'h00260001);
pulp_write32(axi_m, 32'h6600151c, 32'h00260002);
pulp_write32(axi_m, 32'h66001520, 32'h00260003);
pulp_write32(axi_m, 32'h66001524, 32'h00260004);
pulp_write32(axi_m, 32'h66001528, 32'h00260005);
pulp_write32(axi_m, 32'h6600152c, 32'h00260006);
pulp_write32(axi_m, 32'h66001530, 32'h00260007);
pulp_write32(axi_m, 32'h66001534, 32'h00260008);
pulp_write32(axi_m, 32'h66001538, 32'h00260009);
pulp_write32(axi_m, 32'h6600153c, 32'h0026000a);
pulp_write32(axi_m, 32'h66001540, 32'h0026000b);
pulp_write32(axi_m, 32'h66001544, 32'h0026000c);
pulp_write32(axi_m, 32'h66001548, 32'h0026000d);
pulp_write32(axi_m, 32'h6600154c, 32'h0026000e);
pulp_write32(axi_m, 32'h66001550, 32'h0026000f);

pulp_write32(axi_m, 32'h66001554, 32'd39);
pulp_write32(axi_m, 32'h66001558, 32'd1);
pulp_write32(axi_m, 32'h6600155c, 32'h80001a60);
pulp_write32(axi_m, 32'h66001a60, 32'h8000166c);
pulp_write32(axi_m, 32'h660015a0, 32'h00270000);
pulp_write32(axi_m, 32'h660015a4, 32'h00270001);
pulp_write32(axi_m, 32'h660015a8, 32'h00270002);
pulp_write32(axi_m, 32'h660015ac, 32'h00270003);
pulp_write32(axi_m, 32'h660015b0, 32'h00270004);
pulp_write32(axi_m, 32'h660015b4, 32'h00270005);
pulp_write32(axi_m, 32'h660015b8, 32'h00270006);
pulp_write32(axi_m, 32'h660015bc, 32'h00270007);
pulp_write32(axi_m, 32'h660015c0, 32'h00270008);
pulp_write32(axi_m, 32'h660015c4, 32'h00270009);
pulp_write32(axi_m, 32'h660015c8, 32'h0027000a);
pulp_write32(axi_m, 32'h660015cc, 32'h0027000b);
pulp_write32(axi_m, 32'h660015d0, 32'h0027000c);
pulp_write32(axi_m, 32'h660015d4, 32'h0027000d);
pulp_write32(axi_m, 32'h660015d8, 32'h0027000e);
pulp_write32(axi_m, 32'h660015dc, 32'h0027000f);

pulp_write32(axi_m, 32'h660015e0, 32'd40);
pulp_write32(axi_m, 32'h660015e4, 32'd1);
pulp_write32(axi_m, 32'h660015e8, 32'h80001a68);
pulp_write32(axi_m, 32'h66001a68, 32'h8000166c);
pulp_write32(axi_m, 32'h6600162c, 32'h00280000);
pulp_write32(axi_m, 32'h66001630, 32'h00280001);
pulp_write32(axi_m, 32'h66001634, 32'h00280002);
pulp_write32(axi_m, 32'h66001638, 32'h00280003);
pulp_write32(axi_m, 32'h6600163c, 32'h00280004);
pulp_write32(axi_m, 32'h66001640, 32'h00280005);
pulp_write32(axi_m, 32'h66001644, 32'h00280006);
pulp_write32(axi_m, 32'h66001648, 32'h00280007);
pulp_write32(axi_m, 32'h6600164c, 32'h00280008);
pulp_write32(axi_m, 32'h66001650, 32'h00280009);
pulp_write32(axi_m, 32'h66001654, 32'h0028000a);
pulp_write32(axi_m, 32'h66001658, 32'h0028000b);
pulp_write32(axi_m, 32'h6600165c, 32'h0028000c);
pulp_write32(axi_m, 32'h66001660, 32'h0028000d);
pulp_write32(axi_m, 32'h66001664, 32'h0028000e);
pulp_write32(axi_m, 32'h66001668, 32'h0028000f);

pulp_write32(axi_m, 32'h6600166c, 32'd41);
pulp_write32(axi_m, 32'h66001670, 32'd0);
pulp_write32(axi_m, 32'h660016b8, 32'h00290000);
pulp_write32(axi_m, 32'h660016bc, 32'h00290001);
pulp_write32(axi_m, 32'h660016c0, 32'h00290002);
pulp_write32(axi_m, 32'h660016c4, 32'h00290003);
pulp_write32(axi_m, 32'h660016c8, 32'h00290004);
pulp_write32(axi_m, 32'h660016cc, 32'h00290005);
pulp_write32(axi_m, 32'h660016d0, 32'h00290006);
pulp_write32(axi_m, 32'h660016d4, 32'h00290007);
pulp_write32(axi_m, 32'h660016d8, 32'h00290008);
pulp_write32(axi_m, 32'h660016dc, 32'h00290009);
pulp_write32(axi_m, 32'h660016e0, 32'h0029000a);
pulp_write32(axi_m, 32'h660016e4, 32'h0029000b);
pulp_write32(axi_m, 32'h660016e8, 32'h0029000c);
pulp_write32(axi_m, 32'h660016ec, 32'h0029000d);
pulp_write32(axi_m, 32'h660016f0, 32'h0029000e);
pulp_write32(axi_m, 32'h660016f4, 32'h0029000f);

pulp_write32(axi_m, 32'h660016f8, 32'd42);
pulp_write32(axi_m, 32'h660016fc, 32'd1);
pulp_write32(axi_m, 32'h66001700, 32'h80001a70);
pulp_write32(axi_m, 32'h66001a70, 32'h80001784);
pulp_write32(axi_m, 32'h66001744, 32'h002a0000);
pulp_write32(axi_m, 32'h66001748, 32'h002a0001);
pulp_write32(axi_m, 32'h6600174c, 32'h002a0002);
pulp_write32(axi_m, 32'h66001750, 32'h002a0003);
pulp_write32(axi_m, 32'h66001754, 32'h002a0004);
pulp_write32(axi_m, 32'h66001758, 32'h002a0005);
pulp_write32(axi_m, 32'h6600175c, 32'h002a0006);
pulp_write32(axi_m, 32'h66001760, 32'h002a0007);
pulp_write32(axi_m, 32'h66001764, 32'h002a0008);
pulp_write32(axi_m, 32'h66001768, 32'h002a0009);
pulp_write32(axi_m, 32'h6600176c, 32'h002a000a);
pulp_write32(axi_m, 32'h66001770, 32'h002a000b);
pulp_write32(axi_m, 32'h66001774, 32'h002a000c);
pulp_write32(axi_m, 32'h66001778, 32'h002a000d);
pulp_write32(axi_m, 32'h6600177c, 32'h002a000e);
pulp_write32(axi_m, 32'h66001780, 32'h002a000f);

pulp_write32(axi_m, 32'h66001784, 32'd43);
pulp_write32(axi_m, 32'h66001788, 32'd1);
pulp_write32(axi_m, 32'h6600178c, 32'h80001a78);
pulp_write32(axi_m, 32'h66001a78, 32'h8000189c);
pulp_write32(axi_m, 32'h660017d0, 32'h002b0000);
pulp_write32(axi_m, 32'h660017d4, 32'h002b0001);
pulp_write32(axi_m, 32'h660017d8, 32'h002b0002);
pulp_write32(axi_m, 32'h660017dc, 32'h002b0003);
pulp_write32(axi_m, 32'h660017e0, 32'h002b0004);
pulp_write32(axi_m, 32'h660017e4, 32'h002b0005);
pulp_write32(axi_m, 32'h660017e8, 32'h002b0006);
pulp_write32(axi_m, 32'h660017ec, 32'h002b0007);
pulp_write32(axi_m, 32'h660017f0, 32'h002b0008);
pulp_write32(axi_m, 32'h660017f4, 32'h002b0009);
pulp_write32(axi_m, 32'h660017f8, 32'h002b000a);
pulp_write32(axi_m, 32'h660017fc, 32'h002b000b);
pulp_write32(axi_m, 32'h66001800, 32'h002b000c);
pulp_write32(axi_m, 32'h66001804, 32'h002b000d);
pulp_write32(axi_m, 32'h66001808, 32'h002b000e);
pulp_write32(axi_m, 32'h6600180c, 32'h002b000f);

pulp_write32(axi_m, 32'h66001810, 32'd44);
pulp_write32(axi_m, 32'h66001814, 32'd1);
pulp_write32(axi_m, 32'h66001818, 32'h80001a80);
pulp_write32(axi_m, 32'h66001a80, 32'h8000189c);
pulp_write32(axi_m, 32'h6600185c, 32'h002c0000);
pulp_write32(axi_m, 32'h66001860, 32'h002c0001);
pulp_write32(axi_m, 32'h66001864, 32'h002c0002);
pulp_write32(axi_m, 32'h66001868, 32'h002c0003);
pulp_write32(axi_m, 32'h6600186c, 32'h002c0004);
pulp_write32(axi_m, 32'h66001870, 32'h002c0005);
pulp_write32(axi_m, 32'h66001874, 32'h002c0006);
pulp_write32(axi_m, 32'h66001878, 32'h002c0007);
pulp_write32(axi_m, 32'h6600187c, 32'h002c0008);
pulp_write32(axi_m, 32'h66001880, 32'h002c0009);
pulp_write32(axi_m, 32'h66001884, 32'h002c000a);
pulp_write32(axi_m, 32'h66001888, 32'h002c000b);
pulp_write32(axi_m, 32'h6600188c, 32'h002c000c);
pulp_write32(axi_m, 32'h66001890, 32'h002c000d);
pulp_write32(axi_m, 32'h66001894, 32'h002c000e);
pulp_write32(axi_m, 32'h66001898, 32'h002c000f);

pulp_write32(axi_m, 32'h6600189c, 32'd45);
pulp_write32(axi_m, 32'h660018a0, 32'd0);
pulp_write32(axi_m, 32'h660018e8, 32'h002d0000);
pulp_write32(axi_m, 32'h660018ec, 32'h002d0001);
pulp_write32(axi_m, 32'h660018f0, 32'h002d0002);
pulp_write32(axi_m, 32'h660018f4, 32'h002d0003);
pulp_write32(axi_m, 32'h660018f8, 32'h002d0004);
pulp_write32(axi_m, 32'h660018fc, 32'h002d0005);
pulp_write32(axi_m, 32'h66001900, 32'h002d0006);
pulp_write32(axi_m, 32'h66001904, 32'h002d0007);
pulp_write32(axi_m, 32'h66001908, 32'h002d0008);
pulp_write32(axi_m, 32'h6600190c, 32'h002d0009);
pulp_write32(axi_m, 32'h66001910, 32'h002d000a);
pulp_write32(axi_m, 32'h66001914, 32'h002d000b);
pulp_write32(axi_m, 32'h66001918, 32'h002d000c);
pulp_write32(axi_m, 32'h6600191c, 32'h002d000d);
pulp_write32(axi_m, 32'h66001920, 32'h002d000e);
pulp_write32(axi_m, 32'h66001924, 32'h002d000f);

